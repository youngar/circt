// Standard header to adapt well known macros to our needs.
`ifdef RANDOMIZE_REG_INIT
  `define RANDOMIZE
`endif

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM {$random}
`endif

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifdef PRINTF_COND
  `define PRINTF_COND_ (`PRINTF_COND)
`else
  `define PRINTF_COND_ 1
`endif

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifdef STOP_COND
  `define STOP_COND_ (`STOP_COND)
`else
  `define STOP_COND_ 1
`endif

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifdef RANDOMIZE
  `ifdef VERILATOR
    `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
  `else
    `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
  `endif
`else
  `define INIT_RANDOM_PROLOG_
`endif

module T_28314_ext(	// rob.scala:340:30
  input  [4:0] R0_addr,
  input        R0_en, R0_clk,
  input  [4:0] W0_addr,
  input        W0_en, W0_clk,
  input  [4:0] W0_data, W1_addr,
  input        W1_en, W1_clk,
  input  [4:0] W1_data, W2_addr,
  input        W2_en, W2_clk,
  input  [4:0] W2_data,
  output [4:0] R0_data);

  reg [4:0] Memory[0:23];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
    if (W1_en)
      Memory[W1_addr] <= W1_data;
    if (W2_en)
      Memory[W2_addr] <= W2_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 5'bx;	// rob.scala:340:30
endmodule

module row_metadata_has_brorjalr_ext(	// rob.scala:296:38
  input  [4:0] R0_addr,
  input        R0_en, R0_clk,
  input  [4:0] R1_addr,
  input        R1_en, R1_clk,
  input  [4:0] R2_addr,
  input        R2_en, R2_clk,
  input  [4:0] R3_addr,
  input        R3_en, R3_clk,
  input  [4:0] R4_addr,
  input        R4_en, R4_clk,
  input  [4:0] R5_addr,
  input        R5_en, R5_clk,
  input  [4:0] R6_addr,
  input        R6_en, R6_clk,
  input  [4:0] R7_addr,
  input        R7_en, R7_clk,
  input  [4:0] R8_addr,
  input        R8_en, R8_clk,
  input  [4:0] R9_addr,
  input        R9_en, R9_clk,
  input  [4:0] R10_addr,
  input        R10_en, R10_clk,
  input  [4:0] R11_addr,
  input        R11_en, R11_clk,
  input  [4:0] R12_addr,
  input        R12_en, R12_clk,
  input  [4:0] R13_addr,
  input        R13_en, R13_clk,
  input  [4:0] R14_addr,
  input        R14_en, R14_clk,
  input  [4:0] R15_addr,
  input        R15_en, R15_clk,
  input  [4:0] R16_addr,
  input        R16_en, R16_clk,
  input  [4:0] R17_addr,
  input        R17_en, R17_clk,
  input  [4:0] R18_addr,
  input        R18_en, R18_clk,
  input  [4:0] R19_addr,
  input        R19_en, R19_clk,
  input  [4:0] R20_addr,
  input        R20_en, R20_clk,
  input  [4:0] R21_addr,
  input        R21_en, R21_clk,
  input  [4:0] R22_addr,
  input        R22_en, R22_clk,
  input  [4:0] R23_addr,
  input        R23_en, R23_clk,
  input  [4:0] R24_addr,
  input        R24_en, R24_clk,
  input  [4:0] W0_addr,
  input        W0_en, W0_clk, W0_data,
  input  [4:0] W1_addr,
  input        W1_en, W1_clk, W1_data,
  output       R0_data, R1_data, R2_data, R3_data, R4_data, R5_data, R6_data, R7_data,
  output       R8_data, R9_data, R10_data, R11_data, R12_data, R13_data, R14_data,
  output       R15_data, R16_data, R17_data, R18_data, R19_data, R20_data, R21_data,
  output       R22_data, R23_data, R24_data);

  reg Memory[0:23];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
    if (W1_en)
      Memory[W1_addr] <= W1_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 1'bx;	// rob.scala:296:38
  assign R1_data = R1_en ? Memory[R1_addr] : 1'bx;	// rob.scala:296:38
  assign R2_data = R2_en ? Memory[R2_addr] : 1'bx;	// rob.scala:296:38
  assign R3_data = R3_en ? Memory[R3_addr] : 1'bx;	// rob.scala:296:38
  assign R4_data = R4_en ? Memory[R4_addr] : 1'bx;	// rob.scala:296:38
  assign R5_data = R5_en ? Memory[R5_addr] : 1'bx;	// rob.scala:296:38
  assign R6_data = R6_en ? Memory[R6_addr] : 1'bx;	// rob.scala:296:38
  assign R7_data = R7_en ? Memory[R7_addr] : 1'bx;	// rob.scala:296:38
  assign R8_data = R8_en ? Memory[R8_addr] : 1'bx;	// rob.scala:296:38
  assign R9_data = R9_en ? Memory[R9_addr] : 1'bx;	// rob.scala:296:38
  assign R10_data = R10_en ? Memory[R10_addr] : 1'bx;	// rob.scala:296:38
  assign R11_data = R11_en ? Memory[R11_addr] : 1'bx;	// rob.scala:296:38
  assign R12_data = R12_en ? Memory[R12_addr] : 1'bx;	// rob.scala:296:38
  assign R13_data = R13_en ? Memory[R13_addr] : 1'bx;	// rob.scala:296:38
  assign R14_data = R14_en ? Memory[R14_addr] : 1'bx;	// rob.scala:296:38
  assign R15_data = R15_en ? Memory[R15_addr] : 1'bx;	// rob.scala:296:38
  assign R16_data = R16_en ? Memory[R16_addr] : 1'bx;	// rob.scala:296:38
  assign R17_data = R17_en ? Memory[R17_addr] : 1'bx;	// rob.scala:296:38
  assign R18_data = R18_en ? Memory[R18_addr] : 1'bx;	// rob.scala:296:38
  assign R19_data = R19_en ? Memory[R19_addr] : 1'bx;	// rob.scala:296:38
  assign R20_data = R20_en ? Memory[R20_addr] : 1'bx;	// rob.scala:296:38
  assign R21_data = R21_en ? Memory[R21_addr] : 1'bx;	// rob.scala:296:38
  assign R22_data = R22_en ? Memory[R22_addr] : 1'bx;	// rob.scala:296:38
  assign R23_data = R23_en ? Memory[R23_addr] : 1'bx;	// rob.scala:296:38
  assign R24_data = R24_en ? Memory[R24_addr] : 1'bx;	// rob.scala:296:38
endmodule

module T_28311_ext(	// rob.scala:339:30
  input  [4:0] R0_addr,
  input        R0_en, R0_clk,
  input  [4:0] R1_addr,
  input        R1_en, R1_clk,
  input  [4:0] R2_addr,
  input        R2_en, R2_clk,
  input  [4:0] R3_addr,
  input        R3_en, R3_clk,
  input  [4:0] R4_addr,
  input        R4_en, R4_clk,
  input  [4:0] R5_addr,
  input        R5_en, R5_clk,
  input  [4:0] R6_addr,
  input        R6_en, R6_clk,
  input  [4:0] R7_addr,
  input        R7_en, R7_clk,
  input  [4:0] R8_addr,
  input        R8_en, R8_clk,
  input  [4:0] R9_addr,
  input        R9_en, R9_clk,
  input  [4:0] R10_addr,
  input        R10_en, R10_clk,
  input  [4:0] R11_addr,
  input        R11_en, R11_clk,
  input  [4:0] R12_addr,
  input        R12_en, R12_clk,
  input  [4:0] R13_addr,
  input        R13_en, R13_clk,
  input  [4:0] R14_addr,
  input        R14_en, R14_clk,
  input  [4:0] R15_addr,
  input        R15_en, R15_clk,
  input  [4:0] R16_addr,
  input        R16_en, R16_clk,
  input  [4:0] R17_addr,
  input        R17_en, R17_clk,
  input  [4:0] R18_addr,
  input        R18_en, R18_clk,
  input  [4:0] R19_addr,
  input        R19_en, R19_clk,
  input  [4:0] R20_addr,
  input        R20_en, R20_clk,
  input  [4:0] R21_addr,
  input        R21_en, R21_clk,
  input  [4:0] R22_addr,
  input        R22_en, R22_clk,
  input  [4:0] R23_addr,
  input        R23_en, R23_clk,
  input  [4:0] R24_addr,
  input        R24_en, R24_clk,
  input  [4:0] W0_addr,
  input        W0_en, W0_clk, W0_data,
  input  [4:0] W1_addr,
  input        W1_en, W1_clk, W1_data,
  input  [4:0] W2_addr,
  input        W2_en, W2_clk, W2_data,
  input  [4:0] W3_addr,
  input        W3_en, W3_clk, W3_data,
  output       R0_data, R1_data, R2_data, R3_data, R4_data, R5_data, R6_data, R7_data,
  output       R8_data, R9_data, R10_data, R11_data, R12_data, R13_data, R14_data,
  output       R15_data, R16_data, R17_data, R18_data, R19_data, R20_data, R21_data,
  output       R22_data, R23_data, R24_data);

  reg Memory[0:23];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
    if (W1_en)
      Memory[W1_addr] <= W1_data;
    if (W2_en)
      Memory[W2_addr] <= W2_data;
    if (W3_en)
      Memory[W3_addr] <= W3_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 1'bx;	// rob.scala:339:30
  assign R1_data = R1_en ? Memory[R1_addr] : 1'bx;	// rob.scala:339:30
  assign R2_data = R2_en ? Memory[R2_addr] : 1'bx;	// rob.scala:339:30
  assign R3_data = R3_en ? Memory[R3_addr] : 1'bx;	// rob.scala:339:30
  assign R4_data = R4_en ? Memory[R4_addr] : 1'bx;	// rob.scala:339:30
  assign R5_data = R5_en ? Memory[R5_addr] : 1'bx;	// rob.scala:339:30
  assign R6_data = R6_en ? Memory[R6_addr] : 1'bx;	// rob.scala:339:30
  assign R7_data = R7_en ? Memory[R7_addr] : 1'bx;	// rob.scala:339:30
  assign R8_data = R8_en ? Memory[R8_addr] : 1'bx;	// rob.scala:339:30
  assign R9_data = R9_en ? Memory[R9_addr] : 1'bx;	// rob.scala:339:30
  assign R10_data = R10_en ? Memory[R10_addr] : 1'bx;	// rob.scala:339:30
  assign R11_data = R11_en ? Memory[R11_addr] : 1'bx;	// rob.scala:339:30
  assign R12_data = R12_en ? Memory[R12_addr] : 1'bx;	// rob.scala:339:30
  assign R13_data = R13_en ? Memory[R13_addr] : 1'bx;	// rob.scala:339:30
  assign R14_data = R14_en ? Memory[R14_addr] : 1'bx;	// rob.scala:339:30
  assign R15_data = R15_en ? Memory[R15_addr] : 1'bx;	// rob.scala:339:30
  assign R16_data = R16_en ? Memory[R16_addr] : 1'bx;	// rob.scala:339:30
  assign R17_data = R17_en ? Memory[R17_addr] : 1'bx;	// rob.scala:339:30
  assign R18_data = R18_en ? Memory[R18_addr] : 1'bx;	// rob.scala:339:30
  assign R19_data = R19_en ? Memory[R19_addr] : 1'bx;	// rob.scala:339:30
  assign R20_data = R20_en ? Memory[R20_addr] : 1'bx;	// rob.scala:339:30
  assign R21_data = R21_en ? Memory[R21_addr] : 1'bx;	// rob.scala:339:30
  assign R22_data = R22_en ? Memory[R22_addr] : 1'bx;	// rob.scala:339:30
  assign R23_data = R23_en ? Memory[R23_addr] : 1'bx;	// rob.scala:339:30
  assign R24_data = R24_en ? Memory[R24_addr] : 1'bx;	// rob.scala:339:30
endmodule

module T_23710_ext(	// rob.scala:335:30
  input  [4:0] R0_addr,
  input        R0_en, R0_clk,
  input  [4:0] R1_addr,
  input        R1_en, R1_clk,
  input  [4:0] R2_addr,
  input        R2_en, R2_clk,
  input  [4:0] R3_addr,
  input        R3_en, R3_clk,
  input  [4:0] R4_addr,
  input        R4_en, R4_clk,
  input  [4:0] R5_addr,
  input        R5_en, R5_clk,
  input  [4:0] R6_addr,
  input        R6_en, R6_clk,
  input  [4:0] R7_addr,
  input        R7_en, R7_clk,
  input  [4:0] R8_addr,
  input        R8_en, R8_clk,
  input  [4:0] R9_addr,
  input        R9_en, R9_clk,
  input  [4:0] R10_addr,
  input        R10_en, R10_clk,
  input  [4:0] R11_addr,
  input        R11_en, R11_clk,
  input  [4:0] R12_addr,
  input        R12_en, R12_clk,
  input  [4:0] R13_addr,
  input        R13_en, R13_clk,
  input  [4:0] R14_addr,
  input        R14_en, R14_clk,
  input  [4:0] R15_addr,
  input        R15_en, R15_clk,
  input  [4:0] R16_addr,
  input        R16_en, R16_clk,
  input  [4:0] R17_addr,
  input        R17_en, R17_clk,
  input  [4:0] R18_addr,
  input        R18_en, R18_clk,
  input  [4:0] R19_addr,
  input        R19_en, R19_clk,
  input  [4:0] R20_addr,
  input        R20_en, R20_clk,
  input  [4:0] R21_addr,
  input        R21_en, R21_clk,
  input  [4:0] R22_addr,
  input        R22_en, R22_clk,
  input  [4:0] R23_addr,
  input        R23_en, R23_clk,
  input  [4:0] R24_addr,
  input        R24_en, R24_clk,
  input  [4:0] W0_addr,
  input        W0_en, W0_clk, W0_data,
  input  [4:0] W1_addr,
  input        W1_en, W1_clk, W1_data,
  input  [4:0] W2_addr,
  input        W2_en, W2_clk, W2_data,
  input  [4:0] W3_addr,
  input        W3_en, W3_clk, W3_data,
  input  [4:0] W4_addr,
  input        W4_en, W4_clk, W4_data,
  output       R0_data, R1_data, R2_data, R3_data, R4_data, R5_data, R6_data, R7_data,
  output       R8_data, R9_data, R10_data, R11_data, R12_data, R13_data, R14_data,
  output       R15_data, R16_data, R17_data, R18_data, R19_data, R20_data, R21_data,
  output       R22_data, R23_data, R24_data);

  reg Memory[0:23];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
    if (W1_en)
      Memory[W1_addr] <= W1_data;
    if (W2_en)
      Memory[W2_addr] <= W2_data;
    if (W3_en)
      Memory[W3_addr] <= W3_data;
    if (W4_en)
      Memory[W4_addr] <= W4_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 1'bx;	// rob.scala:335:30
  assign R1_data = R1_en ? Memory[R1_addr] : 1'bx;	// rob.scala:335:30
  assign R2_data = R2_en ? Memory[R2_addr] : 1'bx;	// rob.scala:335:30
  assign R3_data = R3_en ? Memory[R3_addr] : 1'bx;	// rob.scala:335:30
  assign R4_data = R4_en ? Memory[R4_addr] : 1'bx;	// rob.scala:335:30
  assign R5_data = R5_en ? Memory[R5_addr] : 1'bx;	// rob.scala:335:30
  assign R6_data = R6_en ? Memory[R6_addr] : 1'bx;	// rob.scala:335:30
  assign R7_data = R7_en ? Memory[R7_addr] : 1'bx;	// rob.scala:335:30
  assign R8_data = R8_en ? Memory[R8_addr] : 1'bx;	// rob.scala:335:30
  assign R9_data = R9_en ? Memory[R9_addr] : 1'bx;	// rob.scala:335:30
  assign R10_data = R10_en ? Memory[R10_addr] : 1'bx;	// rob.scala:335:30
  assign R11_data = R11_en ? Memory[R11_addr] : 1'bx;	// rob.scala:335:30
  assign R12_data = R12_en ? Memory[R12_addr] : 1'bx;	// rob.scala:335:30
  assign R13_data = R13_en ? Memory[R13_addr] : 1'bx;	// rob.scala:335:30
  assign R14_data = R14_en ? Memory[R14_addr] : 1'bx;	// rob.scala:335:30
  assign R15_data = R15_en ? Memory[R15_addr] : 1'bx;	// rob.scala:335:30
  assign R16_data = R16_en ? Memory[R16_addr] : 1'bx;	// rob.scala:335:30
  assign R17_data = R17_en ? Memory[R17_addr] : 1'bx;	// rob.scala:335:30
  assign R18_data = R18_en ? Memory[R18_addr] : 1'bx;	// rob.scala:335:30
  assign R19_data = R19_en ? Memory[R19_addr] : 1'bx;	// rob.scala:335:30
  assign R20_data = R20_en ? Memory[R20_addr] : 1'bx;	// rob.scala:335:30
  assign R21_data = R21_en ? Memory[R21_addr] : 1'bx;	// rob.scala:335:30
  assign R22_data = R22_en ? Memory[R22_addr] : 1'bx;	// rob.scala:335:30
  assign R23_data = R23_en ? Memory[R23_addr] : 1'bx;	// rob.scala:335:30
  assign R24_data = R24_en ? Memory[R24_addr] : 1'bx;	// rob.scala:335:30
endmodule

module row_metadata_brob_idx_ext(	// rob.scala:295:35
  input  [4:0] R0_addr,
  input        R0_en, R0_clk,
  input  [4:0] R1_addr,
  input        R1_en, R1_clk,
  input  [4:0] R2_addr,
  input        R2_en, R2_clk,
  input  [4:0] R3_addr,
  input        R3_en, R3_clk,
  input  [4:0] R4_addr,
  input        R4_en, R4_clk,
  input  [4:0] R5_addr,
  input        R5_en, R5_clk,
  input  [4:0] R6_addr,
  input        R6_en, R6_clk,
  input  [4:0] R7_addr,
  input        R7_en, R7_clk,
  input  [4:0] R8_addr,
  input        R8_en, R8_clk,
  input  [4:0] R9_addr,
  input        R9_en, R9_clk,
  input  [4:0] R10_addr,
  input        R10_en, R10_clk,
  input  [4:0] R11_addr,
  input        R11_en, R11_clk,
  input  [4:0] R12_addr,
  input        R12_en, R12_clk,
  input  [4:0] R13_addr,
  input        R13_en, R13_clk,
  input  [4:0] R14_addr,
  input        R14_en, R14_clk,
  input  [4:0] R15_addr,
  input        R15_en, R15_clk,
  input  [4:0] R16_addr,
  input        R16_en, R16_clk,
  input  [4:0] R17_addr,
  input        R17_en, R17_clk,
  input  [4:0] R18_addr,
  input        R18_en, R18_clk,
  input  [4:0] R19_addr,
  input        R19_en, R19_clk,
  input  [4:0] R20_addr,
  input        R20_en, R20_clk,
  input  [4:0] R21_addr,
  input        R21_en, R21_clk,
  input  [4:0] R22_addr,
  input        R22_en, R22_clk,
  input  [4:0] R23_addr,
  input        R23_en, R23_clk,
  input  [4:0] R24_addr,
  input        R24_en, R24_clk,
  input  [4:0] R25_addr,
  input        R25_en, R25_clk,
  input  [4:0] W0_addr,
  input        W0_en, W0_clk,
  input  [4:0] W0_data,
  output [4:0] R0_data, R1_data, R2_data, R3_data, R4_data, R5_data, R6_data, R7_data,
  output [4:0] R8_data, R9_data, R10_data, R11_data, R12_data, R13_data, R14_data,
  output [4:0] R15_data, R16_data, R17_data, R18_data, R19_data, R20_data, R21_data,
  output [4:0] R22_data, R23_data, R24_data, R25_data);

  reg [4:0] Memory[0:23];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 5'bx;	// rob.scala:295:35
  assign R1_data = R1_en ? Memory[R1_addr] : 5'bx;	// rob.scala:295:35
  assign R2_data = R2_en ? Memory[R2_addr] : 5'bx;	// rob.scala:295:35
  assign R3_data = R3_en ? Memory[R3_addr] : 5'bx;	// rob.scala:295:35
  assign R4_data = R4_en ? Memory[R4_addr] : 5'bx;	// rob.scala:295:35
  assign R5_data = R5_en ? Memory[R5_addr] : 5'bx;	// rob.scala:295:35
  assign R6_data = R6_en ? Memory[R6_addr] : 5'bx;	// rob.scala:295:35
  assign R7_data = R7_en ? Memory[R7_addr] : 5'bx;	// rob.scala:295:35
  assign R8_data = R8_en ? Memory[R8_addr] : 5'bx;	// rob.scala:295:35
  assign R9_data = R9_en ? Memory[R9_addr] : 5'bx;	// rob.scala:295:35
  assign R10_data = R10_en ? Memory[R10_addr] : 5'bx;	// rob.scala:295:35
  assign R11_data = R11_en ? Memory[R11_addr] : 5'bx;	// rob.scala:295:35
  assign R12_data = R12_en ? Memory[R12_addr] : 5'bx;	// rob.scala:295:35
  assign R13_data = R13_en ? Memory[R13_addr] : 5'bx;	// rob.scala:295:35
  assign R14_data = R14_en ? Memory[R14_addr] : 5'bx;	// rob.scala:295:35
  assign R15_data = R15_en ? Memory[R15_addr] : 5'bx;	// rob.scala:295:35
  assign R16_data = R16_en ? Memory[R16_addr] : 5'bx;	// rob.scala:295:35
  assign R17_data = R17_en ? Memory[R17_addr] : 5'bx;	// rob.scala:295:35
  assign R18_data = R18_en ? Memory[R18_addr] : 5'bx;	// rob.scala:295:35
  assign R19_data = R19_en ? Memory[R19_addr] : 5'bx;	// rob.scala:295:35
  assign R20_data = R20_en ? Memory[R20_addr] : 5'bx;	// rob.scala:295:35
  assign R21_data = R21_en ? Memory[R21_addr] : 5'bx;	// rob.scala:295:35
  assign R22_data = R22_en ? Memory[R22_addr] : 5'bx;	// rob.scala:295:35
  assign R23_data = R23_en ? Memory[R23_addr] : 5'bx;	// rob.scala:295:35
  assign R24_data = R24_en ? Memory[R24_addr] : 5'bx;	// rob.scala:295:35
  assign R25_data = R25_en ? Memory[R25_addr] : 5'bx;	// rob.scala:295:35
endmodule

module T_23555_ext(	// rob.scala:894:22
  input  [3:0]  R0_addr,
  input         R0_en, R0_clk,
  input  [3:0]  R1_addr,
  input         R1_en, R1_clk,
  input  [3:0]  R2_addr,
  input         R2_en, R2_clk,
  input  [3:0]  R3_addr,
  input         R3_en, R3_clk,
  input  [3:0]  R4_addr,
  input         R4_en, R4_clk,
  input  [3:0]  R5_addr,
  input         R5_en, R5_clk,
  input  [3:0]  R6_addr,
  input         R6_en, R6_clk,
  input  [3:0]  R7_addr,
  input         R7_en, R7_clk,
  input  [3:0]  R8_addr,
  input         R8_en, R8_clk,
  input  [3:0]  R9_addr,
  input         R9_en, R9_clk,
  input  [3:0]  R10_addr,
  input         R10_en, R10_clk,
  input  [3:0]  R11_addr,
  input         R11_en, R11_clk,
  input  [3:0]  R12_addr,
  input         R12_en, R12_clk,
  input  [3:0]  R13_addr,
  input         R13_en, R13_clk,
  input  [3:0]  R14_addr,
  input         R14_en, R14_clk,
  input  [3:0]  R15_addr,
  input         R15_en, R15_clk,
  input  [3:0]  R16_addr,
  input         R16_en, R16_clk,
  input  [3:0]  R17_addr,
  input         R17_en, R17_clk,
  input  [3:0]  R18_addr,
  input         R18_en, R18_clk,
  input  [3:0]  R19_addr,
  input         R19_en, R19_clk,
  input  [3:0]  R20_addr,
  input         R20_en, R20_clk,
  input  [3:0]  R21_addr,
  input         R21_en, R21_clk,
  input  [3:0]  R22_addr,
  input         R22_en, R22_clk,
  input  [3:0]  R23_addr,
  input         R23_en, R23_clk,
  input  [3:0]  R24_addr,
  input         R24_en, R24_clk,
  input  [3:0]  R25_addr,
  input         R25_en, R25_clk,
  input  [3:0]  R26_addr,
  input         R26_en, R26_clk,
  input  [3:0]  R27_addr,
  input         R27_en, R27_clk,
  input  [3:0]  R28_addr,
  input         R28_en, R28_clk,
  input  [3:0]  R29_addr,
  input         R29_en, R29_clk,
  input  [3:0]  R30_addr,
  input         R30_en, R30_clk,
  input  [3:0]  R31_addr,
  input         R31_en, R31_clk,
  input  [3:0]  R32_addr,
  input         R32_en, R32_clk,
  input  [3:0]  R33_addr,
  input         R33_en, R33_clk,
  input  [3:0]  R34_addr,
  input         R34_en, R34_clk,
  input  [3:0]  R35_addr,
  input         R35_en, R35_clk,
  input  [3:0]  R36_addr,
  input         R36_en, R36_clk,
  input  [3:0]  R37_addr,
  input         R37_en, R37_clk,
  input  [3:0]  R38_addr,
  input         R38_en, R38_clk,
  input  [3:0]  R39_addr,
  input         R39_en, R39_clk,
  input  [3:0]  R40_addr,
  input         R40_en, R40_clk,
  input  [3:0]  R41_addr,
  input         R41_en, R41_clk,
  input  [3:0]  R42_addr,
  input         R42_en, R42_clk,
  input  [3:0]  R43_addr,
  input         R43_en, R43_clk,
  input  [3:0]  R44_addr,
  input         R44_en, R44_clk,
  input  [3:0]  R45_addr,
  input         R45_en, R45_clk,
  input  [3:0]  R46_addr,
  input         R46_en, R46_clk,
  input  [3:0]  R47_addr,
  input         R47_en, R47_clk,
  input  [3:0]  R48_addr,
  input         R48_en, R48_clk,
  input  [3:0]  R49_addr,
  input         R49_en, R49_clk,
  input  [3:0]  W0_addr,
  input         W0_en, W0_clk,
  input  [36:0] W0_data,
  output [36:0] R0_data, R1_data, R2_data, R3_data, R4_data, R5_data, R6_data, R7_data,
  output [36:0] R8_data, R9_data, R10_data, R11_data, R12_data, R13_data, R14_data,
  output [36:0] R15_data, R16_data, R17_data, R18_data, R19_data, R20_data, R21_data,
  output [36:0] R22_data, R23_data, R24_data, R25_data, R26_data, R27_data, R28_data,
  output [36:0] R29_data, R30_data, R31_data, R32_data, R33_data, R34_data, R35_data,
  output [36:0] R36_data, R37_data, R38_data, R39_data, R40_data, R41_data, R42_data,
  output [36:0] R43_data, R44_data, R45_data, R46_data, R47_data, R48_data, R49_data);

  reg [36:0] Memory[0:11];

  always @(posedge W0_clk) begin
    if (W0_en)
      Memory[W0_addr] <= W0_data;
  end // always @(posedge)
  assign R0_data = R0_en ? Memory[R0_addr] : 37'bx;	// rob.scala:894:22
  assign R1_data = R1_en ? Memory[R1_addr] : 37'bx;	// rob.scala:894:22
  assign R2_data = R2_en ? Memory[R2_addr] : 37'bx;	// rob.scala:894:22
  assign R3_data = R3_en ? Memory[R3_addr] : 37'bx;	// rob.scala:894:22
  assign R4_data = R4_en ? Memory[R4_addr] : 37'bx;	// rob.scala:894:22
  assign R5_data = R5_en ? Memory[R5_addr] : 37'bx;	// rob.scala:894:22
  assign R6_data = R6_en ? Memory[R6_addr] : 37'bx;	// rob.scala:894:22
  assign R7_data = R7_en ? Memory[R7_addr] : 37'bx;	// rob.scala:894:22
  assign R8_data = R8_en ? Memory[R8_addr] : 37'bx;	// rob.scala:894:22
  assign R9_data = R9_en ? Memory[R9_addr] : 37'bx;	// rob.scala:894:22
  assign R10_data = R10_en ? Memory[R10_addr] : 37'bx;	// rob.scala:894:22
  assign R11_data = R11_en ? Memory[R11_addr] : 37'bx;	// rob.scala:894:22
  assign R12_data = R12_en ? Memory[R12_addr] : 37'bx;	// rob.scala:894:22
  assign R13_data = R13_en ? Memory[R13_addr] : 37'bx;	// rob.scala:894:22
  assign R14_data = R14_en ? Memory[R14_addr] : 37'bx;	// rob.scala:894:22
  assign R15_data = R15_en ? Memory[R15_addr] : 37'bx;	// rob.scala:894:22
  assign R16_data = R16_en ? Memory[R16_addr] : 37'bx;	// rob.scala:894:22
  assign R17_data = R17_en ? Memory[R17_addr] : 37'bx;	// rob.scala:894:22
  assign R18_data = R18_en ? Memory[R18_addr] : 37'bx;	// rob.scala:894:22
  assign R19_data = R19_en ? Memory[R19_addr] : 37'bx;	// rob.scala:894:22
  assign R20_data = R20_en ? Memory[R20_addr] : 37'bx;	// rob.scala:894:22
  assign R21_data = R21_en ? Memory[R21_addr] : 37'bx;	// rob.scala:894:22
  assign R22_data = R22_en ? Memory[R22_addr] : 37'bx;	// rob.scala:894:22
  assign R23_data = R23_en ? Memory[R23_addr] : 37'bx;	// rob.scala:894:22
  assign R24_data = R24_en ? Memory[R24_addr] : 37'bx;	// rob.scala:894:22
  assign R25_data = R25_en ? Memory[R25_addr] : 37'bx;	// rob.scala:894:22
  assign R26_data = R26_en ? Memory[R26_addr] : 37'bx;	// rob.scala:894:22
  assign R27_data = R27_en ? Memory[R27_addr] : 37'bx;	// rob.scala:894:22
  assign R28_data = R28_en ? Memory[R28_addr] : 37'bx;	// rob.scala:894:22
  assign R29_data = R29_en ? Memory[R29_addr] : 37'bx;	// rob.scala:894:22
  assign R30_data = R30_en ? Memory[R30_addr] : 37'bx;	// rob.scala:894:22
  assign R31_data = R31_en ? Memory[R31_addr] : 37'bx;	// rob.scala:894:22
  assign R32_data = R32_en ? Memory[R32_addr] : 37'bx;	// rob.scala:894:22
  assign R33_data = R33_en ? Memory[R33_addr] : 37'bx;	// rob.scala:894:22
  assign R34_data = R34_en ? Memory[R34_addr] : 37'bx;	// rob.scala:894:22
  assign R35_data = R35_en ? Memory[R35_addr] : 37'bx;	// rob.scala:894:22
  assign R36_data = R36_en ? Memory[R36_addr] : 37'bx;	// rob.scala:894:22
  assign R37_data = R37_en ? Memory[R37_addr] : 37'bx;	// rob.scala:894:22
  assign R38_data = R38_en ? Memory[R38_addr] : 37'bx;	// rob.scala:894:22
  assign R39_data = R39_en ? Memory[R39_addr] : 37'bx;	// rob.scala:894:22
  assign R40_data = R40_en ? Memory[R40_addr] : 37'bx;	// rob.scala:894:22
  assign R41_data = R41_en ? Memory[R41_addr] : 37'bx;	// rob.scala:894:22
  assign R42_data = R42_en ? Memory[R42_addr] : 37'bx;	// rob.scala:894:22
  assign R43_data = R43_en ? Memory[R43_addr] : 37'bx;	// rob.scala:894:22
  assign R44_data = R44_en ? Memory[R44_addr] : 37'bx;	// rob.scala:894:22
  assign R45_data = R45_en ? Memory[R45_addr] : 37'bx;	// rob.scala:894:22
  assign R46_data = R46_en ? Memory[R46_addr] : 37'bx;	// rob.scala:894:22
  assign R47_data = R47_en ? Memory[R47_addr] : 37'bx;	// rob.scala:894:22
  assign R48_data = R48_en ? Memory[R48_addr] : 37'bx;	// rob.scala:894:22
  assign R49_data = R49_en ? Memory[R49_addr] : 37'bx;	// rob.scala:894:22
endmodule

module Rob(	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  input         clk, reset, io_dis_valids_0, io_dis_valids_1, io_dis_uops_0_valid,
  input  [1:0]  io_dis_uops_0_iw_state,
  input  [8:0]  io_dis_uops_0_uopc,
  input  [31:0] io_dis_uops_0_inst,
  input  [39:0] io_dis_uops_0_pc,
  input  [7:0]  io_dis_uops_0_fu_code,
  input  [3:0]  io_dis_uops_0_ctrl_br_type,
  input  [1:0]  io_dis_uops_0_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_0_ctrl_op2_sel, io_dis_uops_0_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_0_ctrl_op_fcn,
  input         io_dis_uops_0_ctrl_fcn_dw, io_dis_uops_0_ctrl_rf_wen,
  input  [2:0]  io_dis_uops_0_ctrl_csr_cmd,
  input         io_dis_uops_0_ctrl_is_load, io_dis_uops_0_ctrl_is_sta,
  input         io_dis_uops_0_ctrl_is_std,
  input  [1:0]  io_dis_uops_0_wakeup_delay,
  input         io_dis_uops_0_allocate_brtag, io_dis_uops_0_is_br_or_jmp,
  input         io_dis_uops_0_is_jump, io_dis_uops_0_is_jal, io_dis_uops_0_is_ret,
  input         io_dis_uops_0_is_call,
  input  [7:0]  io_dis_uops_0_br_mask,
  input  [2:0]  io_dis_uops_0_br_tag,
  input         io_dis_uops_0_br_prediction_bpd_predict_val,
  input         io_dis_uops_0_br_prediction_bpd_predict_taken,
  input         io_dis_uops_0_br_prediction_btb_hit,
  input         io_dis_uops_0_br_prediction_btb_predicted,
  input         io_dis_uops_0_br_prediction_is_br_or_jalr,
  input         io_dis_uops_0_stat_brjmp_mispredicted, io_dis_uops_0_stat_btb_made_pred,
  input         io_dis_uops_0_stat_btb_mispredicted, io_dis_uops_0_stat_bpd_made_pred,
  input         io_dis_uops_0_stat_bpd_mispredicted,
  input  [2:0]  io_dis_uops_0_fetch_pc_lob,
  input  [19:0] io_dis_uops_0_imm_packed,
  input  [11:0] io_dis_uops_0_csr_addr,
  input  [5:0]  io_dis_uops_0_rob_idx,
  input  [3:0]  io_dis_uops_0_ldq_idx, io_dis_uops_0_stq_idx,
  input  [4:0]  io_dis_uops_0_brob_idx,
  input  [6:0]  io_dis_uops_0_pdst, io_dis_uops_0_pop1, io_dis_uops_0_pop2,
  input  [6:0]  io_dis_uops_0_pop3,
  input         io_dis_uops_0_prs1_busy, io_dis_uops_0_prs2_busy,
  input         io_dis_uops_0_prs3_busy,
  input  [6:0]  io_dis_uops_0_stale_pdst,
  input         io_dis_uops_0_exception,
  input  [63:0] io_dis_uops_0_exc_cause,
  input         io_dis_uops_0_bypassable,
  input  [3:0]  io_dis_uops_0_mem_cmd,
  input  [2:0]  io_dis_uops_0_mem_typ,
  input         io_dis_uops_0_is_fence, io_dis_uops_0_is_fencei, io_dis_uops_0_is_store,
  input         io_dis_uops_0_is_amo, io_dis_uops_0_is_load, io_dis_uops_0_is_unique,
  input         io_dis_uops_0_flush_on_commit,
  input  [5:0]  io_dis_uops_0_ldst, io_dis_uops_0_lrs1, io_dis_uops_0_lrs2,
  input  [5:0]  io_dis_uops_0_lrs3,
  input         io_dis_uops_0_ldst_val,
  input  [1:0]  io_dis_uops_0_dst_rtype, io_dis_uops_0_lrs1_rtype,
  input  [1:0]  io_dis_uops_0_lrs2_rtype,
  input         io_dis_uops_0_frs3_en, io_dis_uops_0_fp_val, io_dis_uops_0_fp_single,
  input         io_dis_uops_0_xcpt_if, io_dis_uops_0_replay_if,
  input  [63:0] io_dis_uops_0_debug_wdata,
  input  [31:0] io_dis_uops_0_debug_events_fetch_seq,
  input         io_dis_uops_1_valid,
  input  [1:0]  io_dis_uops_1_iw_state,
  input  [8:0]  io_dis_uops_1_uopc,
  input  [31:0] io_dis_uops_1_inst,
  input  [39:0] io_dis_uops_1_pc,
  input  [7:0]  io_dis_uops_1_fu_code,
  input  [3:0]  io_dis_uops_1_ctrl_br_type,
  input  [1:0]  io_dis_uops_1_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_1_ctrl_op2_sel, io_dis_uops_1_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_1_ctrl_op_fcn,
  input         io_dis_uops_1_ctrl_fcn_dw, io_dis_uops_1_ctrl_rf_wen,
  input  [2:0]  io_dis_uops_1_ctrl_csr_cmd,
  input         io_dis_uops_1_ctrl_is_load, io_dis_uops_1_ctrl_is_sta,
  input         io_dis_uops_1_ctrl_is_std,
  input  [1:0]  io_dis_uops_1_wakeup_delay,
  input         io_dis_uops_1_allocate_brtag, io_dis_uops_1_is_br_or_jmp,
  input         io_dis_uops_1_is_jump, io_dis_uops_1_is_jal, io_dis_uops_1_is_ret,
  input         io_dis_uops_1_is_call,
  input  [7:0]  io_dis_uops_1_br_mask,
  input  [2:0]  io_dis_uops_1_br_tag,
  input         io_dis_uops_1_br_prediction_bpd_predict_val,
  input         io_dis_uops_1_br_prediction_bpd_predict_taken,
  input         io_dis_uops_1_br_prediction_btb_hit,
  input         io_dis_uops_1_br_prediction_btb_predicted,
  input         io_dis_uops_1_br_prediction_is_br_or_jalr,
  input         io_dis_uops_1_stat_brjmp_mispredicted, io_dis_uops_1_stat_btb_made_pred,
  input         io_dis_uops_1_stat_btb_mispredicted, io_dis_uops_1_stat_bpd_made_pred,
  input         io_dis_uops_1_stat_bpd_mispredicted,
  input  [2:0]  io_dis_uops_1_fetch_pc_lob,
  input  [19:0] io_dis_uops_1_imm_packed,
  input  [11:0] io_dis_uops_1_csr_addr,
  input  [5:0]  io_dis_uops_1_rob_idx,
  input  [3:0]  io_dis_uops_1_ldq_idx, io_dis_uops_1_stq_idx,
  input  [4:0]  io_dis_uops_1_brob_idx,
  input  [6:0]  io_dis_uops_1_pdst, io_dis_uops_1_pop1, io_dis_uops_1_pop2,
  input  [6:0]  io_dis_uops_1_pop3,
  input         io_dis_uops_1_prs1_busy, io_dis_uops_1_prs2_busy,
  input         io_dis_uops_1_prs3_busy,
  input  [6:0]  io_dis_uops_1_stale_pdst,
  input         io_dis_uops_1_exception,
  input  [63:0] io_dis_uops_1_exc_cause,
  input         io_dis_uops_1_bypassable,
  input  [3:0]  io_dis_uops_1_mem_cmd,
  input  [2:0]  io_dis_uops_1_mem_typ,
  input         io_dis_uops_1_is_fence, io_dis_uops_1_is_fencei, io_dis_uops_1_is_store,
  input         io_dis_uops_1_is_amo, io_dis_uops_1_is_load, io_dis_uops_1_is_unique,
  input         io_dis_uops_1_flush_on_commit,
  input  [5:0]  io_dis_uops_1_ldst, io_dis_uops_1_lrs1, io_dis_uops_1_lrs2,
  input  [5:0]  io_dis_uops_1_lrs3,
  input         io_dis_uops_1_ldst_val,
  input  [1:0]  io_dis_uops_1_dst_rtype, io_dis_uops_1_lrs1_rtype,
  input  [1:0]  io_dis_uops_1_lrs2_rtype,
  input         io_dis_uops_1_frs3_en, io_dis_uops_1_fp_val, io_dis_uops_1_fp_single,
  input         io_dis_uops_1_xcpt_if, io_dis_uops_1_replay_if,
  input  [63:0] io_dis_uops_1_debug_wdata,
  input  [31:0] io_dis_uops_1_debug_events_fetch_seq,
  input         io_dis_has_br_or_jalr_in_packet, io_dis_partial_stall, io_dis_new_packet,
  input         io_wb_resps_0_valid, io_wb_resps_0_bits_uop_valid,
  input  [1:0]  io_wb_resps_0_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_0_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_uop_inst,
  input  [39:0] io_wb_resps_0_bits_uop_pc,
  input  [7:0]  io_wb_resps_0_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_op2_sel, io_wb_resps_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_uop_ctrl_fcn_dw, io_wb_resps_0_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_0_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_uop_ctrl_is_load, io_wb_resps_0_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_uop_wakeup_delay,
  input         io_wb_resps_0_bits_uop_allocate_brtag,
  input         io_wb_resps_0_bits_uop_is_br_or_jmp, io_wb_resps_0_bits_uop_is_jump,
  input         io_wb_resps_0_bits_uop_is_jal, io_wb_resps_0_bits_uop_is_ret,
  input         io_wb_resps_0_bits_uop_is_call,
  input  [7:0]  io_wb_resps_0_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_uop_br_tag,
  input         io_wb_resps_0_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_0_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_0_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_0_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_0_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_0_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_0_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_0_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_0_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_0_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_0_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_0_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_0_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_0_bits_uop_ldq_idx, io_wb_resps_0_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_0_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_0_bits_uop_pdst, io_wb_resps_0_bits_uop_pop1,
  input  [6:0]  io_wb_resps_0_bits_uop_pop2, io_wb_resps_0_bits_uop_pop3,
  input         io_wb_resps_0_bits_uop_prs1_busy, io_wb_resps_0_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_0_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_0_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_0_bits_uop_mem_typ,
  input         io_wb_resps_0_bits_uop_is_fence, io_wb_resps_0_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_uop_is_store, io_wb_resps_0_bits_uop_is_amo,
  input         io_wb_resps_0_bits_uop_is_load, io_wb_resps_0_bits_uop_is_unique,
  input         io_wb_resps_0_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_0_bits_uop_ldst, io_wb_resps_0_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_uop_lrs2, io_wb_resps_0_bits_uop_lrs3,
  input         io_wb_resps_0_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_uop_dst_rtype, io_wb_resps_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_uop_frs3_en, io_wb_resps_0_bits_uop_fp_val,
  input         io_wb_resps_0_bits_uop_fp_single, io_wb_resps_0_bits_uop_xcpt_if,
  input         io_wb_resps_0_bits_uop_replay_if,
  input  [63:0] io_wb_resps_0_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_0_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_0_bits_data,
  input         io_wb_resps_0_bits_fflags_valid,
  input         io_wb_resps_0_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_0_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_0_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_0_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_0_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_0_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_0_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_0_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_0_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_0_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_0_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_0_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_0_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_0_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_0_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_0_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_0_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_0_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_0_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_0_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_0_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_0_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_0_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_0_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_0_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_0_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_0_bits_fflags_bits_flags,
  input         io_wb_resps_1_valid, io_wb_resps_1_bits_uop_valid,
  input  [1:0]  io_wb_resps_1_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_1_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_uop_inst,
  input  [39:0] io_wb_resps_1_bits_uop_pc,
  input  [7:0]  io_wb_resps_1_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_op2_sel, io_wb_resps_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_uop_ctrl_fcn_dw, io_wb_resps_1_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_1_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_uop_ctrl_is_load, io_wb_resps_1_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_uop_wakeup_delay,
  input         io_wb_resps_1_bits_uop_allocate_brtag,
  input         io_wb_resps_1_bits_uop_is_br_or_jmp, io_wb_resps_1_bits_uop_is_jump,
  input         io_wb_resps_1_bits_uop_is_jal, io_wb_resps_1_bits_uop_is_ret,
  input         io_wb_resps_1_bits_uop_is_call,
  input  [7:0]  io_wb_resps_1_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_uop_br_tag,
  input         io_wb_resps_1_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_1_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_1_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_1_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_1_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_1_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_1_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_1_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_1_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_1_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_1_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_1_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_1_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_1_bits_uop_ldq_idx, io_wb_resps_1_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_1_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_1_bits_uop_pdst, io_wb_resps_1_bits_uop_pop1,
  input  [6:0]  io_wb_resps_1_bits_uop_pop2, io_wb_resps_1_bits_uop_pop3,
  input         io_wb_resps_1_bits_uop_prs1_busy, io_wb_resps_1_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_1_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_1_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_1_bits_uop_mem_typ,
  input         io_wb_resps_1_bits_uop_is_fence, io_wb_resps_1_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_uop_is_store, io_wb_resps_1_bits_uop_is_amo,
  input         io_wb_resps_1_bits_uop_is_load, io_wb_resps_1_bits_uop_is_unique,
  input         io_wb_resps_1_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_1_bits_uop_ldst, io_wb_resps_1_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_uop_lrs2, io_wb_resps_1_bits_uop_lrs3,
  input         io_wb_resps_1_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_uop_dst_rtype, io_wb_resps_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_uop_frs3_en, io_wb_resps_1_bits_uop_fp_val,
  input         io_wb_resps_1_bits_uop_fp_single, io_wb_resps_1_bits_uop_xcpt_if,
  input         io_wb_resps_1_bits_uop_replay_if,
  input  [63:0] io_wb_resps_1_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_1_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_1_bits_data,
  input         io_wb_resps_1_bits_fflags_valid,
  input         io_wb_resps_1_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_1_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_1_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_1_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_1_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_1_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_1_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_1_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_1_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_1_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_1_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_1_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_1_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_1_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_1_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_1_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_1_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_1_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_1_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_1_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_1_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_1_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_1_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_1_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_1_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_1_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_1_bits_fflags_bits_flags,
  input         io_wb_resps_2_valid, io_wb_resps_2_bits_uop_valid,
  input  [1:0]  io_wb_resps_2_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_2_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_uop_inst,
  input  [39:0] io_wb_resps_2_bits_uop_pc,
  input  [7:0]  io_wb_resps_2_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_op2_sel, io_wb_resps_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_uop_ctrl_fcn_dw, io_wb_resps_2_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_2_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_uop_ctrl_is_load, io_wb_resps_2_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_uop_wakeup_delay,
  input         io_wb_resps_2_bits_uop_allocate_brtag,
  input         io_wb_resps_2_bits_uop_is_br_or_jmp, io_wb_resps_2_bits_uop_is_jump,
  input         io_wb_resps_2_bits_uop_is_jal, io_wb_resps_2_bits_uop_is_ret,
  input         io_wb_resps_2_bits_uop_is_call,
  input  [7:0]  io_wb_resps_2_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_uop_br_tag,
  input         io_wb_resps_2_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_2_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_2_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_2_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_2_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_2_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_2_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_2_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_2_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_2_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_2_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_2_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_2_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_2_bits_uop_ldq_idx, io_wb_resps_2_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_2_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_2_bits_uop_pdst, io_wb_resps_2_bits_uop_pop1,
  input  [6:0]  io_wb_resps_2_bits_uop_pop2, io_wb_resps_2_bits_uop_pop3,
  input         io_wb_resps_2_bits_uop_prs1_busy, io_wb_resps_2_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_2_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_2_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_2_bits_uop_mem_typ,
  input         io_wb_resps_2_bits_uop_is_fence, io_wb_resps_2_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_uop_is_store, io_wb_resps_2_bits_uop_is_amo,
  input         io_wb_resps_2_bits_uop_is_load, io_wb_resps_2_bits_uop_is_unique,
  input         io_wb_resps_2_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_2_bits_uop_ldst, io_wb_resps_2_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_uop_lrs2, io_wb_resps_2_bits_uop_lrs3,
  input         io_wb_resps_2_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_uop_dst_rtype, io_wb_resps_2_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_uop_frs3_en, io_wb_resps_2_bits_uop_fp_val,
  input         io_wb_resps_2_bits_uop_fp_single, io_wb_resps_2_bits_uop_xcpt_if,
  input         io_wb_resps_2_bits_uop_replay_if,
  input  [63:0] io_wb_resps_2_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_2_bits_uop_debug_events_fetch_seq,
  input  [64:0] io_wb_resps_2_bits_data,
  input         io_wb_resps_2_bits_fflags_valid,
  input         io_wb_resps_2_bits_fflags_bits_uop_valid,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_iw_state,
  input  [8:0]  io_wb_resps_2_bits_fflags_bits_uop_uopc,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_inst,
  input  [39:0] io_wb_resps_2_bits_fflags_bits_uop_pc,
  input  [7:0]  io_wb_resps_2_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_fcn_dw,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_load,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_wb_resps_2_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_wakeup_delay,
  input         io_wb_resps_2_bits_fflags_bits_uop_allocate_brtag,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_br_or_jmp,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jump,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_jal,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_ret,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_call,
  input  [7:0]  io_wb_resps_2_bits_fflags_bits_uop_br_mask,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_br_tag,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_bpd_predict_val,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_bpd_predict_taken,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_btb_hit,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_btb_predicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_br_prediction_is_br_or_jalr,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_brjmp_mispredicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_btb_made_pred,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_btb_mispredicted,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_bpd_made_pred,
  input         io_wb_resps_2_bits_fflags_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_fetch_pc_lob,
  input  [19:0] io_wb_resps_2_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_wb_resps_2_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_rob_idx,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_ldq_idx,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_stq_idx,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_uop_brob_idx,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop1,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop2,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_pop3,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs1_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs2_busy,
  input         io_wb_resps_2_bits_fflags_bits_uop_prs3_busy,
  input  [6:0]  io_wb_resps_2_bits_fflags_bits_uop_stale_pdst,
  input         io_wb_resps_2_bits_fflags_bits_uop_exception,
  input  [63:0] io_wb_resps_2_bits_fflags_bits_uop_exc_cause,
  input         io_wb_resps_2_bits_fflags_bits_uop_bypassable,
  input  [3:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_cmd,
  input  [2:0]  io_wb_resps_2_bits_fflags_bits_uop_mem_typ,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fence,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_fencei,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_store,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_amo,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_load,
  input         io_wb_resps_2_bits_fflags_bits_uop_is_unique,
  input         io_wb_resps_2_bits_fflags_bits_uop_flush_on_commit,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs3,
  input         io_wb_resps_2_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_wb_resps_2_bits_fflags_bits_uop_lrs2_rtype,
  input         io_wb_resps_2_bits_fflags_bits_uop_frs3_en,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_val,
  input         io_wb_resps_2_bits_fflags_bits_uop_fp_single,
  input         io_wb_resps_2_bits_fflags_bits_uop_xcpt_if,
  input         io_wb_resps_2_bits_fflags_bits_uop_replay_if,
  input  [63:0] io_wb_resps_2_bits_fflags_bits_uop_debug_wdata,
  input  [31:0] io_wb_resps_2_bits_fflags_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_wb_resps_2_bits_fflags_bits_flags,
  input         io_debug_wb_valids_0, io_debug_wb_valids_1, io_debug_wb_valids_2,
  input  [63:0] io_debug_wb_wdata_0, io_debug_wb_wdata_1, io_debug_wb_wdata_2,
  input         io_fflags_0_valid, io_fflags_0_bits_uop_valid,
  input  [1:0]  io_fflags_0_bits_uop_iw_state,
  input  [8:0]  io_fflags_0_bits_uop_uopc,
  input  [31:0] io_fflags_0_bits_uop_inst,
  input  [39:0] io_fflags_0_bits_uop_pc,
  input  [7:0]  io_fflags_0_bits_uop_fu_code,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_op2_sel, io_fflags_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_0_bits_uop_ctrl_op_fcn,
  input         io_fflags_0_bits_uop_ctrl_fcn_dw, io_fflags_0_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_fflags_0_bits_uop_ctrl_csr_cmd,
  input         io_fflags_0_bits_uop_ctrl_is_load, io_fflags_0_bits_uop_ctrl_is_sta,
  input         io_fflags_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_0_bits_uop_wakeup_delay,
  input         io_fflags_0_bits_uop_allocate_brtag, io_fflags_0_bits_uop_is_br_or_jmp,
  input         io_fflags_0_bits_uop_is_jump, io_fflags_0_bits_uop_is_jal,
  input         io_fflags_0_bits_uop_is_ret, io_fflags_0_bits_uop_is_call,
  input  [7:0]  io_fflags_0_bits_uop_br_mask,
  input  [2:0]  io_fflags_0_bits_uop_br_tag,
  input         io_fflags_0_bits_uop_br_prediction_bpd_predict_val,
  input         io_fflags_0_bits_uop_br_prediction_bpd_predict_taken,
  input         io_fflags_0_bits_uop_br_prediction_btb_hit,
  input         io_fflags_0_bits_uop_br_prediction_btb_predicted,
  input         io_fflags_0_bits_uop_br_prediction_is_br_or_jalr,
  input         io_fflags_0_bits_uop_stat_brjmp_mispredicted,
  input         io_fflags_0_bits_uop_stat_btb_made_pred,
  input         io_fflags_0_bits_uop_stat_btb_mispredicted,
  input         io_fflags_0_bits_uop_stat_bpd_made_pred,
  input         io_fflags_0_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_fflags_0_bits_uop_fetch_pc_lob,
  input  [19:0] io_fflags_0_bits_uop_imm_packed,
  input  [11:0] io_fflags_0_bits_uop_csr_addr,
  input  [5:0]  io_fflags_0_bits_uop_rob_idx,
  input  [3:0]  io_fflags_0_bits_uop_ldq_idx, io_fflags_0_bits_uop_stq_idx,
  input  [4:0]  io_fflags_0_bits_uop_brob_idx,
  input  [6:0]  io_fflags_0_bits_uop_pdst, io_fflags_0_bits_uop_pop1,
  input  [6:0]  io_fflags_0_bits_uop_pop2, io_fflags_0_bits_uop_pop3,
  input         io_fflags_0_bits_uop_prs1_busy, io_fflags_0_bits_uop_prs2_busy,
  input         io_fflags_0_bits_uop_prs3_busy,
  input  [6:0]  io_fflags_0_bits_uop_stale_pdst,
  input         io_fflags_0_bits_uop_exception,
  input  [63:0] io_fflags_0_bits_uop_exc_cause,
  input         io_fflags_0_bits_uop_bypassable,
  input  [3:0]  io_fflags_0_bits_uop_mem_cmd,
  input  [2:0]  io_fflags_0_bits_uop_mem_typ,
  input         io_fflags_0_bits_uop_is_fence, io_fflags_0_bits_uop_is_fencei,
  input         io_fflags_0_bits_uop_is_store, io_fflags_0_bits_uop_is_amo,
  input         io_fflags_0_bits_uop_is_load, io_fflags_0_bits_uop_is_unique,
  input         io_fflags_0_bits_uop_flush_on_commit,
  input  [5:0]  io_fflags_0_bits_uop_ldst, io_fflags_0_bits_uop_lrs1,
  input  [5:0]  io_fflags_0_bits_uop_lrs2, io_fflags_0_bits_uop_lrs3,
  input         io_fflags_0_bits_uop_ldst_val,
  input  [1:0]  io_fflags_0_bits_uop_dst_rtype, io_fflags_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_0_bits_uop_lrs2_rtype,
  input         io_fflags_0_bits_uop_frs3_en, io_fflags_0_bits_uop_fp_val,
  input         io_fflags_0_bits_uop_fp_single, io_fflags_0_bits_uop_xcpt_if,
  input         io_fflags_0_bits_uop_replay_if,
  input  [63:0] io_fflags_0_bits_uop_debug_wdata,
  input  [31:0] io_fflags_0_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_1_valid, io_fflags_1_bits_uop_valid,
  input  [1:0]  io_fflags_1_bits_uop_iw_state,
  input  [8:0]  io_fflags_1_bits_uop_uopc,
  input  [31:0] io_fflags_1_bits_uop_inst,
  input  [39:0] io_fflags_1_bits_uop_pc,
  input  [7:0]  io_fflags_1_bits_uop_fu_code,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_fflags_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_op2_sel, io_fflags_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_fflags_1_bits_uop_ctrl_op_fcn,
  input         io_fflags_1_bits_uop_ctrl_fcn_dw, io_fflags_1_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_fflags_1_bits_uop_ctrl_csr_cmd,
  input         io_fflags_1_bits_uop_ctrl_is_load, io_fflags_1_bits_uop_ctrl_is_sta,
  input         io_fflags_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_fflags_1_bits_uop_wakeup_delay,
  input         io_fflags_1_bits_uop_allocate_brtag, io_fflags_1_bits_uop_is_br_or_jmp,
  input         io_fflags_1_bits_uop_is_jump, io_fflags_1_bits_uop_is_jal,
  input         io_fflags_1_bits_uop_is_ret, io_fflags_1_bits_uop_is_call,
  input  [7:0]  io_fflags_1_bits_uop_br_mask,
  input  [2:0]  io_fflags_1_bits_uop_br_tag,
  input         io_fflags_1_bits_uop_br_prediction_bpd_predict_val,
  input         io_fflags_1_bits_uop_br_prediction_bpd_predict_taken,
  input         io_fflags_1_bits_uop_br_prediction_btb_hit,
  input         io_fflags_1_bits_uop_br_prediction_btb_predicted,
  input         io_fflags_1_bits_uop_br_prediction_is_br_or_jalr,
  input         io_fflags_1_bits_uop_stat_brjmp_mispredicted,
  input         io_fflags_1_bits_uop_stat_btb_made_pred,
  input         io_fflags_1_bits_uop_stat_btb_mispredicted,
  input         io_fflags_1_bits_uop_stat_bpd_made_pred,
  input         io_fflags_1_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_fflags_1_bits_uop_fetch_pc_lob,
  input  [19:0] io_fflags_1_bits_uop_imm_packed,
  input  [11:0] io_fflags_1_bits_uop_csr_addr,
  input  [5:0]  io_fflags_1_bits_uop_rob_idx,
  input  [3:0]  io_fflags_1_bits_uop_ldq_idx, io_fflags_1_bits_uop_stq_idx,
  input  [4:0]  io_fflags_1_bits_uop_brob_idx,
  input  [6:0]  io_fflags_1_bits_uop_pdst, io_fflags_1_bits_uop_pop1,
  input  [6:0]  io_fflags_1_bits_uop_pop2, io_fflags_1_bits_uop_pop3,
  input         io_fflags_1_bits_uop_prs1_busy, io_fflags_1_bits_uop_prs2_busy,
  input         io_fflags_1_bits_uop_prs3_busy,
  input  [6:0]  io_fflags_1_bits_uop_stale_pdst,
  input         io_fflags_1_bits_uop_exception,
  input  [63:0] io_fflags_1_bits_uop_exc_cause,
  input         io_fflags_1_bits_uop_bypassable,
  input  [3:0]  io_fflags_1_bits_uop_mem_cmd,
  input  [2:0]  io_fflags_1_bits_uop_mem_typ,
  input         io_fflags_1_bits_uop_is_fence, io_fflags_1_bits_uop_is_fencei,
  input         io_fflags_1_bits_uop_is_store, io_fflags_1_bits_uop_is_amo,
  input         io_fflags_1_bits_uop_is_load, io_fflags_1_bits_uop_is_unique,
  input         io_fflags_1_bits_uop_flush_on_commit,
  input  [5:0]  io_fflags_1_bits_uop_ldst, io_fflags_1_bits_uop_lrs1,
  input  [5:0]  io_fflags_1_bits_uop_lrs2, io_fflags_1_bits_uop_lrs3,
  input         io_fflags_1_bits_uop_ldst_val,
  input  [1:0]  io_fflags_1_bits_uop_dst_rtype, io_fflags_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_fflags_1_bits_uop_lrs2_rtype,
  input         io_fflags_1_bits_uop_frs3_en, io_fflags_1_bits_uop_fp_val,
  input         io_fflags_1_bits_uop_fp_single, io_fflags_1_bits_uop_xcpt_if,
  input         io_fflags_1_bits_uop_replay_if,
  input  [63:0] io_fflags_1_bits_uop_debug_wdata,
  input  [31:0] io_fflags_1_bits_uop_debug_events_fetch_seq,
  input  [4:0]  io_fflags_1_bits_flags,
  input         io_lxcpt_valid, io_lxcpt_bits_uop_valid,
  input  [1:0]  io_lxcpt_bits_uop_iw_state,
  input  [8:0]  io_lxcpt_bits_uop_uopc,
  input  [31:0] io_lxcpt_bits_uop_inst,
  input  [39:0] io_lxcpt_bits_uop_pc,
  input  [7:0]  io_lxcpt_bits_uop_fu_code,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_lxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_op2_sel, io_lxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_lxcpt_bits_uop_ctrl_op_fcn,
  input         io_lxcpt_bits_uop_ctrl_fcn_dw, io_lxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_lxcpt_bits_uop_ctrl_csr_cmd,
  input         io_lxcpt_bits_uop_ctrl_is_load, io_lxcpt_bits_uop_ctrl_is_sta,
  input         io_lxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_lxcpt_bits_uop_wakeup_delay,
  input         io_lxcpt_bits_uop_allocate_brtag, io_lxcpt_bits_uop_is_br_or_jmp,
  input         io_lxcpt_bits_uop_is_jump, io_lxcpt_bits_uop_is_jal,
  input         io_lxcpt_bits_uop_is_ret, io_lxcpt_bits_uop_is_call,
  input  [7:0]  io_lxcpt_bits_uop_br_mask,
  input  [2:0]  io_lxcpt_bits_uop_br_tag,
  input         io_lxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_lxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_lxcpt_bits_uop_br_prediction_btb_hit,
  input         io_lxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_lxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_lxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_lxcpt_bits_uop_stat_btb_made_pred,
  input         io_lxcpt_bits_uop_stat_btb_mispredicted,
  input         io_lxcpt_bits_uop_stat_bpd_made_pred,
  input         io_lxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_lxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_lxcpt_bits_uop_imm_packed,
  input  [11:0] io_lxcpt_bits_uop_csr_addr,
  input  [5:0]  io_lxcpt_bits_uop_rob_idx,
  input  [3:0]  io_lxcpt_bits_uop_ldq_idx, io_lxcpt_bits_uop_stq_idx,
  input  [4:0]  io_lxcpt_bits_uop_brob_idx,
  input  [6:0]  io_lxcpt_bits_uop_pdst, io_lxcpt_bits_uop_pop1, io_lxcpt_bits_uop_pop2,
  input  [6:0]  io_lxcpt_bits_uop_pop3,
  input         io_lxcpt_bits_uop_prs1_busy, io_lxcpt_bits_uop_prs2_busy,
  input         io_lxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_lxcpt_bits_uop_stale_pdst,
  input         io_lxcpt_bits_uop_exception,
  input  [63:0] io_lxcpt_bits_uop_exc_cause,
  input         io_lxcpt_bits_uop_bypassable,
  input  [3:0]  io_lxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_lxcpt_bits_uop_mem_typ,
  input         io_lxcpt_bits_uop_is_fence, io_lxcpt_bits_uop_is_fencei,
  input         io_lxcpt_bits_uop_is_store, io_lxcpt_bits_uop_is_amo,
  input         io_lxcpt_bits_uop_is_load, io_lxcpt_bits_uop_is_unique,
  input         io_lxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_lxcpt_bits_uop_ldst, io_lxcpt_bits_uop_lrs1, io_lxcpt_bits_uop_lrs2,
  input  [5:0]  io_lxcpt_bits_uop_lrs3,
  input         io_lxcpt_bits_uop_ldst_val,
  input  [1:0]  io_lxcpt_bits_uop_dst_rtype, io_lxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_lxcpt_bits_uop_lrs2_rtype,
  input         io_lxcpt_bits_uop_frs3_en, io_lxcpt_bits_uop_fp_val,
  input         io_lxcpt_bits_uop_fp_single, io_lxcpt_bits_uop_xcpt_if,
  input         io_lxcpt_bits_uop_replay_if,
  input  [63:0] io_lxcpt_bits_uop_debug_wdata,
  input  [31:0] io_lxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_bxcpt_valid, io_bxcpt_bits_uop_valid,
  input  [1:0]  io_bxcpt_bits_uop_iw_state,
  input  [8:0]  io_bxcpt_bits_uop_uopc,
  input  [31:0] io_bxcpt_bits_uop_inst,
  input  [39:0] io_bxcpt_bits_uop_pc,
  input  [7:0]  io_bxcpt_bits_uop_fu_code,
  input  [3:0]  io_bxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_bxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bxcpt_bits_uop_ctrl_op2_sel, io_bxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bxcpt_bits_uop_ctrl_op_fcn,
  input         io_bxcpt_bits_uop_ctrl_fcn_dw, io_bxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_bxcpt_bits_uop_ctrl_csr_cmd,
  input         io_bxcpt_bits_uop_ctrl_is_load, io_bxcpt_bits_uop_ctrl_is_sta,
  input         io_bxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_bxcpt_bits_uop_wakeup_delay,
  input         io_bxcpt_bits_uop_allocate_brtag, io_bxcpt_bits_uop_is_br_or_jmp,
  input         io_bxcpt_bits_uop_is_jump, io_bxcpt_bits_uop_is_jal,
  input         io_bxcpt_bits_uop_is_ret, io_bxcpt_bits_uop_is_call,
  input  [7:0]  io_bxcpt_bits_uop_br_mask,
  input  [2:0]  io_bxcpt_bits_uop_br_tag,
  input         io_bxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_bxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_bxcpt_bits_uop_br_prediction_btb_hit,
  input         io_bxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_bxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_bxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_bxcpt_bits_uop_stat_btb_made_pred,
  input         io_bxcpt_bits_uop_stat_btb_mispredicted,
  input         io_bxcpt_bits_uop_stat_bpd_made_pred,
  input         io_bxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_bxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_bxcpt_bits_uop_imm_packed,
  input  [11:0] io_bxcpt_bits_uop_csr_addr,
  input  [5:0]  io_bxcpt_bits_uop_rob_idx,
  input  [3:0]  io_bxcpt_bits_uop_ldq_idx, io_bxcpt_bits_uop_stq_idx,
  input  [4:0]  io_bxcpt_bits_uop_brob_idx,
  input  [6:0]  io_bxcpt_bits_uop_pdst, io_bxcpt_bits_uop_pop1, io_bxcpt_bits_uop_pop2,
  input  [6:0]  io_bxcpt_bits_uop_pop3,
  input         io_bxcpt_bits_uop_prs1_busy, io_bxcpt_bits_uop_prs2_busy,
  input         io_bxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_bxcpt_bits_uop_stale_pdst,
  input         io_bxcpt_bits_uop_exception,
  input  [63:0] io_bxcpt_bits_uop_exc_cause,
  input         io_bxcpt_bits_uop_bypassable,
  input  [3:0]  io_bxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_bxcpt_bits_uop_mem_typ,
  input         io_bxcpt_bits_uop_is_fence, io_bxcpt_bits_uop_is_fencei,
  input         io_bxcpt_bits_uop_is_store, io_bxcpt_bits_uop_is_amo,
  input         io_bxcpt_bits_uop_is_load, io_bxcpt_bits_uop_is_unique,
  input         io_bxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_bxcpt_bits_uop_ldst, io_bxcpt_bits_uop_lrs1, io_bxcpt_bits_uop_lrs2,
  input  [5:0]  io_bxcpt_bits_uop_lrs3,
  input         io_bxcpt_bits_uop_ldst_val,
  input  [1:0]  io_bxcpt_bits_uop_dst_rtype, io_bxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_bxcpt_bits_uop_lrs2_rtype,
  input         io_bxcpt_bits_uop_frs3_en, io_bxcpt_bits_uop_fp_val,
  input         io_bxcpt_bits_uop_fp_single, io_bxcpt_bits_uop_xcpt_if,
  input         io_bxcpt_bits_uop_replay_if,
  input  [63:0] io_bxcpt_bits_uop_debug_wdata,
  input  [31:0] io_bxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_bxcpt_bits_cause,
  input  [39:0] io_bxcpt_bits_badvaddr,
  input         io_cxcpt_valid, io_cxcpt_bits_uop_valid,
  input  [1:0]  io_cxcpt_bits_uop_iw_state,
  input  [8:0]  io_cxcpt_bits_uop_uopc,
  input  [31:0] io_cxcpt_bits_uop_inst,
  input  [39:0] io_cxcpt_bits_uop_pc,
  input  [7:0]  io_cxcpt_bits_uop_fu_code,
  input  [3:0]  io_cxcpt_bits_uop_ctrl_br_type,
  input  [1:0]  io_cxcpt_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_cxcpt_bits_uop_ctrl_op2_sel, io_cxcpt_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_cxcpt_bits_uop_ctrl_op_fcn,
  input         io_cxcpt_bits_uop_ctrl_fcn_dw, io_cxcpt_bits_uop_ctrl_rf_wen,
  input  [2:0]  io_cxcpt_bits_uop_ctrl_csr_cmd,
  input         io_cxcpt_bits_uop_ctrl_is_load, io_cxcpt_bits_uop_ctrl_is_sta,
  input         io_cxcpt_bits_uop_ctrl_is_std,
  input  [1:0]  io_cxcpt_bits_uop_wakeup_delay,
  input         io_cxcpt_bits_uop_allocate_brtag, io_cxcpt_bits_uop_is_br_or_jmp,
  input         io_cxcpt_bits_uop_is_jump, io_cxcpt_bits_uop_is_jal,
  input         io_cxcpt_bits_uop_is_ret, io_cxcpt_bits_uop_is_call,
  input  [7:0]  io_cxcpt_bits_uop_br_mask,
  input  [2:0]  io_cxcpt_bits_uop_br_tag,
  input         io_cxcpt_bits_uop_br_prediction_bpd_predict_val,
  input         io_cxcpt_bits_uop_br_prediction_bpd_predict_taken,
  input         io_cxcpt_bits_uop_br_prediction_btb_hit,
  input         io_cxcpt_bits_uop_br_prediction_btb_predicted,
  input         io_cxcpt_bits_uop_br_prediction_is_br_or_jalr,
  input         io_cxcpt_bits_uop_stat_brjmp_mispredicted,
  input         io_cxcpt_bits_uop_stat_btb_made_pred,
  input         io_cxcpt_bits_uop_stat_btb_mispredicted,
  input         io_cxcpt_bits_uop_stat_bpd_made_pred,
  input         io_cxcpt_bits_uop_stat_bpd_mispredicted,
  input  [2:0]  io_cxcpt_bits_uop_fetch_pc_lob,
  input  [19:0] io_cxcpt_bits_uop_imm_packed,
  input  [11:0] io_cxcpt_bits_uop_csr_addr,
  input  [5:0]  io_cxcpt_bits_uop_rob_idx,
  input  [3:0]  io_cxcpt_bits_uop_ldq_idx, io_cxcpt_bits_uop_stq_idx,
  input  [4:0]  io_cxcpt_bits_uop_brob_idx,
  input  [6:0]  io_cxcpt_bits_uop_pdst, io_cxcpt_bits_uop_pop1, io_cxcpt_bits_uop_pop2,
  input  [6:0]  io_cxcpt_bits_uop_pop3,
  input         io_cxcpt_bits_uop_prs1_busy, io_cxcpt_bits_uop_prs2_busy,
  input         io_cxcpt_bits_uop_prs3_busy,
  input  [6:0]  io_cxcpt_bits_uop_stale_pdst,
  input         io_cxcpt_bits_uop_exception,
  input  [63:0] io_cxcpt_bits_uop_exc_cause,
  input         io_cxcpt_bits_uop_bypassable,
  input  [3:0]  io_cxcpt_bits_uop_mem_cmd,
  input  [2:0]  io_cxcpt_bits_uop_mem_typ,
  input         io_cxcpt_bits_uop_is_fence, io_cxcpt_bits_uop_is_fencei,
  input         io_cxcpt_bits_uop_is_store, io_cxcpt_bits_uop_is_amo,
  input         io_cxcpt_bits_uop_is_load, io_cxcpt_bits_uop_is_unique,
  input         io_cxcpt_bits_uop_flush_on_commit,
  input  [5:0]  io_cxcpt_bits_uop_ldst, io_cxcpt_bits_uop_lrs1, io_cxcpt_bits_uop_lrs2,
  input  [5:0]  io_cxcpt_bits_uop_lrs3,
  input         io_cxcpt_bits_uop_ldst_val,
  input  [1:0]  io_cxcpt_bits_uop_dst_rtype, io_cxcpt_bits_uop_lrs1_rtype,
  input  [1:0]  io_cxcpt_bits_uop_lrs2_rtype,
  input         io_cxcpt_bits_uop_frs3_en, io_cxcpt_bits_uop_fp_val,
  input         io_cxcpt_bits_uop_fp_single, io_cxcpt_bits_uop_xcpt_if,
  input         io_cxcpt_bits_uop_replay_if,
  input  [63:0] io_cxcpt_bits_uop_debug_wdata,
  input  [31:0] io_cxcpt_bits_uop_debug_events_fetch_seq,
  input  [3:0]  io_cxcpt_bits_cause,
  input  [39:0] io_cxcpt_bits_badvaddr,
  input         io_lsu_clr_bsy_valid,
  input  [5:0]  io_lsu_clr_bsy_rob_idx,
  input         io_brinfo_valid, io_brinfo_mispredict,
  input  [7:0]  io_brinfo_mask,
  input  [2:0]  io_brinfo_tag,
  input  [7:0]  io_brinfo_exe_mask,
  input  [5:0]  io_brinfo_rob_idx,
  input  [3:0]  io_brinfo_ldq_idx, io_brinfo_stq_idx,
  input         io_brinfo_taken, io_brinfo_is_jr, io_brinfo_btb_made_pred,
  input         io_brinfo_btb_mispredict, io_brinfo_bpd_made_pred,
  input         io_brinfo_bpd_mispredict,
  input  [5:0]  io_get_pc_rob_idx,
  input  [63:0] io_debug_tsc,
  output [5:0]  io_curr_rob_tail,
  output        io_com_valids_0, io_com_valids_1, io_com_uops_0_valid,
  output [1:0]  io_com_uops_0_iw_state,
  output [8:0]  io_com_uops_0_uopc,
  output [31:0] io_com_uops_0_inst,
  output [39:0] io_com_uops_0_pc,
  output [7:0]  io_com_uops_0_fu_code,
  output [3:0]  io_com_uops_0_ctrl_br_type,
  output [1:0]  io_com_uops_0_ctrl_op1_sel,
  output [2:0]  io_com_uops_0_ctrl_op2_sel, io_com_uops_0_ctrl_imm_sel,
  output [3:0]  io_com_uops_0_ctrl_op_fcn,
  output        io_com_uops_0_ctrl_fcn_dw, io_com_uops_0_ctrl_rf_wen,
  output [2:0]  io_com_uops_0_ctrl_csr_cmd,
  output        io_com_uops_0_ctrl_is_load, io_com_uops_0_ctrl_is_sta,
  output        io_com_uops_0_ctrl_is_std,
  output [1:0]  io_com_uops_0_wakeup_delay,
  output        io_com_uops_0_allocate_brtag, io_com_uops_0_is_br_or_jmp,
  output        io_com_uops_0_is_jump, io_com_uops_0_is_jal, io_com_uops_0_is_ret,
  output        io_com_uops_0_is_call,
  output [7:0]  io_com_uops_0_br_mask,
  output [2:0]  io_com_uops_0_br_tag,
  output        io_com_uops_0_br_prediction_bpd_predict_val,
  output        io_com_uops_0_br_prediction_bpd_predict_taken,
  output        io_com_uops_0_br_prediction_btb_hit,
  output        io_com_uops_0_br_prediction_btb_predicted,
  output        io_com_uops_0_br_prediction_is_br_or_jalr,
  output        io_com_uops_0_stat_brjmp_mispredicted, io_com_uops_0_stat_btb_made_pred,
  output        io_com_uops_0_stat_btb_mispredicted, io_com_uops_0_stat_bpd_made_pred,
  output        io_com_uops_0_stat_bpd_mispredicted,
  output [2:0]  io_com_uops_0_fetch_pc_lob,
  output [19:0] io_com_uops_0_imm_packed,
  output [11:0] io_com_uops_0_csr_addr,
  output [5:0]  io_com_uops_0_rob_idx,
  output [3:0]  io_com_uops_0_ldq_idx, io_com_uops_0_stq_idx,
  output [4:0]  io_com_uops_0_brob_idx,
  output [6:0]  io_com_uops_0_pdst, io_com_uops_0_pop1, io_com_uops_0_pop2,
  output [6:0]  io_com_uops_0_pop3,
  output        io_com_uops_0_prs1_busy, io_com_uops_0_prs2_busy,
  output        io_com_uops_0_prs3_busy,
  output [6:0]  io_com_uops_0_stale_pdst,
  output        io_com_uops_0_exception,
  output [63:0] io_com_uops_0_exc_cause,
  output        io_com_uops_0_bypassable,
  output [3:0]  io_com_uops_0_mem_cmd,
  output [2:0]  io_com_uops_0_mem_typ,
  output        io_com_uops_0_is_fence, io_com_uops_0_is_fencei, io_com_uops_0_is_store,
  output        io_com_uops_0_is_amo, io_com_uops_0_is_load, io_com_uops_0_is_unique,
  output        io_com_uops_0_flush_on_commit,
  output [5:0]  io_com_uops_0_ldst, io_com_uops_0_lrs1, io_com_uops_0_lrs2,
  output [5:0]  io_com_uops_0_lrs3,
  output        io_com_uops_0_ldst_val,
  output [1:0]  io_com_uops_0_dst_rtype, io_com_uops_0_lrs1_rtype,
  output [1:0]  io_com_uops_0_lrs2_rtype,
  output        io_com_uops_0_frs3_en, io_com_uops_0_fp_val, io_com_uops_0_fp_single,
  output        io_com_uops_0_xcpt_if, io_com_uops_0_replay_if,
  output [63:0] io_com_uops_0_debug_wdata,
  output [31:0] io_com_uops_0_debug_events_fetch_seq,
  output        io_com_uops_1_valid,
  output [1:0]  io_com_uops_1_iw_state,
  output [8:0]  io_com_uops_1_uopc,
  output [31:0] io_com_uops_1_inst,
  output [39:0] io_com_uops_1_pc,
  output [7:0]  io_com_uops_1_fu_code,
  output [3:0]  io_com_uops_1_ctrl_br_type,
  output [1:0]  io_com_uops_1_ctrl_op1_sel,
  output [2:0]  io_com_uops_1_ctrl_op2_sel, io_com_uops_1_ctrl_imm_sel,
  output [3:0]  io_com_uops_1_ctrl_op_fcn,
  output        io_com_uops_1_ctrl_fcn_dw, io_com_uops_1_ctrl_rf_wen,
  output [2:0]  io_com_uops_1_ctrl_csr_cmd,
  output        io_com_uops_1_ctrl_is_load, io_com_uops_1_ctrl_is_sta,
  output        io_com_uops_1_ctrl_is_std,
  output [1:0]  io_com_uops_1_wakeup_delay,
  output        io_com_uops_1_allocate_brtag, io_com_uops_1_is_br_or_jmp,
  output        io_com_uops_1_is_jump, io_com_uops_1_is_jal, io_com_uops_1_is_ret,
  output        io_com_uops_1_is_call,
  output [7:0]  io_com_uops_1_br_mask,
  output [2:0]  io_com_uops_1_br_tag,
  output        io_com_uops_1_br_prediction_bpd_predict_val,
  output        io_com_uops_1_br_prediction_bpd_predict_taken,
  output        io_com_uops_1_br_prediction_btb_hit,
  output        io_com_uops_1_br_prediction_btb_predicted,
  output        io_com_uops_1_br_prediction_is_br_or_jalr,
  output        io_com_uops_1_stat_brjmp_mispredicted, io_com_uops_1_stat_btb_made_pred,
  output        io_com_uops_1_stat_btb_mispredicted, io_com_uops_1_stat_bpd_made_pred,
  output        io_com_uops_1_stat_bpd_mispredicted,
  output [2:0]  io_com_uops_1_fetch_pc_lob,
  output [19:0] io_com_uops_1_imm_packed,
  output [11:0] io_com_uops_1_csr_addr,
  output [5:0]  io_com_uops_1_rob_idx,
  output [3:0]  io_com_uops_1_ldq_idx, io_com_uops_1_stq_idx,
  output [4:0]  io_com_uops_1_brob_idx,
  output [6:0]  io_com_uops_1_pdst, io_com_uops_1_pop1, io_com_uops_1_pop2,
  output [6:0]  io_com_uops_1_pop3,
  output        io_com_uops_1_prs1_busy, io_com_uops_1_prs2_busy,
  output        io_com_uops_1_prs3_busy,
  output [6:0]  io_com_uops_1_stale_pdst,
  output        io_com_uops_1_exception,
  output [63:0] io_com_uops_1_exc_cause,
  output        io_com_uops_1_bypassable,
  output [3:0]  io_com_uops_1_mem_cmd,
  output [2:0]  io_com_uops_1_mem_typ,
  output        io_com_uops_1_is_fence, io_com_uops_1_is_fencei, io_com_uops_1_is_store,
  output        io_com_uops_1_is_amo, io_com_uops_1_is_load, io_com_uops_1_is_unique,
  output        io_com_uops_1_flush_on_commit,
  output [5:0]  io_com_uops_1_ldst, io_com_uops_1_lrs1, io_com_uops_1_lrs2,
  output [5:0]  io_com_uops_1_lrs3,
  output        io_com_uops_1_ldst_val,
  output [1:0]  io_com_uops_1_dst_rtype, io_com_uops_1_lrs1_rtype,
  output [1:0]  io_com_uops_1_lrs2_rtype,
  output        io_com_uops_1_frs3_en, io_com_uops_1_fp_val, io_com_uops_1_fp_single,
  output        io_com_uops_1_xcpt_if, io_com_uops_1_replay_if,
  output [63:0] io_com_uops_1_debug_wdata,
  output [31:0] io_com_uops_1_debug_events_fetch_seq,
  output        io_com_fflags_val,
  output [4:0]  io_com_fflags,
  output        io_com_st_mask_0, io_com_st_mask_1, io_com_ld_mask_0, io_com_ld_mask_1,
  output        io_com_load_is_at_rob_head, io_com_exception,
  output [63:0] io_com_exc_cause,
  output        io_com_handling_exc, io_com_rbk_valids_0, io_com_rbk_valids_1,
  output [63:0] io_com_badvaddr,
  output [39:0] io_get_pc_curr_pc,
  output [4:0]  io_get_pc_curr_brob_idx,
  output        io_get_pc_next_val,
  output [39:0] io_get_pc_next_pc,
  output        io_lsu_misspec, io_flush_take_pc,
  output [39:0] io_flush_pc,
  output        io_flush_pipeline, io_flush_brob, io_empty, io_ready,
  output        io_brob_deallocate_valid,
  output [4:0]  io_brob_deallocate_bits_brob_idx,
  output [1:0]  io_debug_state,
  output [5:0]  io_debug_rob_head,
  output        io_debug_xcpt_val, io_debug_xcpt_uop_valid,
  output [1:0]  io_debug_xcpt_uop_iw_state,
  output [8:0]  io_debug_xcpt_uop_uopc,
  output [31:0] io_debug_xcpt_uop_inst,
  output [39:0] io_debug_xcpt_uop_pc,
  output [7:0]  io_debug_xcpt_uop_fu_code,
  output [3:0]  io_debug_xcpt_uop_ctrl_br_type,
  output [1:0]  io_debug_xcpt_uop_ctrl_op1_sel,
  output [2:0]  io_debug_xcpt_uop_ctrl_op2_sel, io_debug_xcpt_uop_ctrl_imm_sel,
  output [3:0]  io_debug_xcpt_uop_ctrl_op_fcn,
  output        io_debug_xcpt_uop_ctrl_fcn_dw, io_debug_xcpt_uop_ctrl_rf_wen,
  output [2:0]  io_debug_xcpt_uop_ctrl_csr_cmd,
  output        io_debug_xcpt_uop_ctrl_is_load, io_debug_xcpt_uop_ctrl_is_sta,
  output        io_debug_xcpt_uop_ctrl_is_std,
  output [1:0]  io_debug_xcpt_uop_wakeup_delay,
  output        io_debug_xcpt_uop_allocate_brtag, io_debug_xcpt_uop_is_br_or_jmp,
  output        io_debug_xcpt_uop_is_jump, io_debug_xcpt_uop_is_jal,
  output        io_debug_xcpt_uop_is_ret, io_debug_xcpt_uop_is_call,
  output [7:0]  io_debug_xcpt_uop_br_mask,
  output [2:0]  io_debug_xcpt_uop_br_tag,
  output        io_debug_xcpt_uop_br_prediction_bpd_predict_val,
  output        io_debug_xcpt_uop_br_prediction_bpd_predict_taken,
  output        io_debug_xcpt_uop_br_prediction_btb_hit,
  output        io_debug_xcpt_uop_br_prediction_btb_predicted,
  output        io_debug_xcpt_uop_br_prediction_is_br_or_jalr,
  output        io_debug_xcpt_uop_stat_brjmp_mispredicted,
  output        io_debug_xcpt_uop_stat_btb_made_pred,
  output        io_debug_xcpt_uop_stat_btb_mispredicted,
  output        io_debug_xcpt_uop_stat_bpd_made_pred,
  output        io_debug_xcpt_uop_stat_bpd_mispredicted,
  output [2:0]  io_debug_xcpt_uop_fetch_pc_lob,
  output [19:0] io_debug_xcpt_uop_imm_packed,
  output [11:0] io_debug_xcpt_uop_csr_addr,
  output [5:0]  io_debug_xcpt_uop_rob_idx,
  output [3:0]  io_debug_xcpt_uop_ldq_idx, io_debug_xcpt_uop_stq_idx,
  output [4:0]  io_debug_xcpt_uop_brob_idx,
  output [6:0]  io_debug_xcpt_uop_pdst, io_debug_xcpt_uop_pop1, io_debug_xcpt_uop_pop2,
  output [6:0]  io_debug_xcpt_uop_pop3,
  output        io_debug_xcpt_uop_prs1_busy, io_debug_xcpt_uop_prs2_busy,
  output        io_debug_xcpt_uop_prs3_busy,
  output [6:0]  io_debug_xcpt_uop_stale_pdst,
  output        io_debug_xcpt_uop_exception,
  output [63:0] io_debug_xcpt_uop_exc_cause,
  output        io_debug_xcpt_uop_bypassable,
  output [3:0]  io_debug_xcpt_uop_mem_cmd,
  output [2:0]  io_debug_xcpt_uop_mem_typ,
  output        io_debug_xcpt_uop_is_fence, io_debug_xcpt_uop_is_fencei,
  output        io_debug_xcpt_uop_is_store, io_debug_xcpt_uop_is_amo,
  output        io_debug_xcpt_uop_is_load, io_debug_xcpt_uop_is_unique,
  output        io_debug_xcpt_uop_flush_on_commit,
  output [5:0]  io_debug_xcpt_uop_ldst, io_debug_xcpt_uop_lrs1, io_debug_xcpt_uop_lrs2,
  output [5:0]  io_debug_xcpt_uop_lrs3,
  output        io_debug_xcpt_uop_ldst_val,
  output [1:0]  io_debug_xcpt_uop_dst_rtype, io_debug_xcpt_uop_lrs1_rtype,
  output [1:0]  io_debug_xcpt_uop_lrs2_rtype,
  output        io_debug_xcpt_uop_frs3_en, io_debug_xcpt_uop_fp_val,
  output        io_debug_xcpt_uop_fp_single, io_debug_xcpt_uop_xcpt_if,
  output        io_debug_xcpt_uop_replay_if,
  output [63:0] io_debug_xcpt_uop_debug_wdata,
  output [31:0] io_debug_xcpt_uop_debug_events_fetch_seq,
  output [63:0] io_debug_xcpt_badvaddr);

  wire        _T;	// rob.scala:716:89
  wire        _T_0;	// rob.scala:509:28
  wire        _T_1;	// rob.scala:509:28
  wire [4:0]  T_40242_R0_data;	// rob.scala:340:30
  wire        T_40239_R0_data;	// rob.scala:339:30
  wire        T_40239_R1_data;	// rob.scala:339:30
  wire        T_40239_R2_data;	// rob.scala:339:30
  wire        T_40239_R3_data;	// rob.scala:339:30
  wire        T_40239_R4_data;	// rob.scala:339:30
  wire        T_40239_R5_data;	// rob.scala:339:30
  wire        T_40239_R6_data;	// rob.scala:339:30
  wire        T_40239_R7_data;	// rob.scala:339:30
  wire        T_40239_R8_data;	// rob.scala:339:30
  wire        T_40239_R9_data;	// rob.scala:339:30
  wire        T_40239_R10_data;	// rob.scala:339:30
  wire        T_40239_R11_data;	// rob.scala:339:30
  wire        T_40239_R12_data;	// rob.scala:339:30
  wire        T_40239_R13_data;	// rob.scala:339:30
  wire        T_40239_R14_data;	// rob.scala:339:30
  wire        T_40239_R15_data;	// rob.scala:339:30
  wire        T_40239_R16_data;	// rob.scala:339:30
  wire        T_40239_R17_data;	// rob.scala:339:30
  wire        T_40239_R18_data;	// rob.scala:339:30
  wire        T_40239_R19_data;	// rob.scala:339:30
  wire        T_40239_R20_data;	// rob.scala:339:30
  wire        T_40239_R21_data;	// rob.scala:339:30
  wire        T_40239_R22_data;	// rob.scala:339:30
  wire        T_40239_R23_data;	// rob.scala:339:30
  wire        T_40239_R24_data;	// rob.scala:339:30
  wire        T_35638_R0_data;	// rob.scala:335:30
  wire        T_35638_R1_data;	// rob.scala:335:30
  wire        T_35638_R2_data;	// rob.scala:335:30
  wire        T_35638_R3_data;	// rob.scala:335:30
  wire        T_35638_R4_data;	// rob.scala:335:30
  wire        T_35638_R5_data;	// rob.scala:335:30
  wire        T_35638_R6_data;	// rob.scala:335:30
  wire        T_35638_R7_data;	// rob.scala:335:30
  wire        T_35638_R8_data;	// rob.scala:335:30
  wire        T_35638_R9_data;	// rob.scala:335:30
  wire        T_35638_R10_data;	// rob.scala:335:30
  wire        T_35638_R11_data;	// rob.scala:335:30
  wire        T_35638_R12_data;	// rob.scala:335:30
  wire        T_35638_R13_data;	// rob.scala:335:30
  wire        T_35638_R14_data;	// rob.scala:335:30
  wire        T_35638_R15_data;	// rob.scala:335:30
  wire        T_35638_R16_data;	// rob.scala:335:30
  wire        T_35638_R17_data;	// rob.scala:335:30
  wire        T_35638_R18_data;	// rob.scala:335:30
  wire        T_35638_R19_data;	// rob.scala:335:30
  wire        T_35638_R20_data;	// rob.scala:335:30
  wire        T_35638_R21_data;	// rob.scala:335:30
  wire        T_35638_R22_data;	// rob.scala:335:30
  wire        T_35638_R23_data;	// rob.scala:335:30
  wire        T_35638_R24_data;	// rob.scala:335:30
  wire [4:0]  T_28314_R0_data;	// rob.scala:340:30
  wire        T_28311_R0_data;	// rob.scala:339:30
  wire        T_28311_R1_data;	// rob.scala:339:30
  wire        T_28311_R2_data;	// rob.scala:339:30
  wire        T_28311_R3_data;	// rob.scala:339:30
  wire        T_28311_R4_data;	// rob.scala:339:30
  wire        T_28311_R5_data;	// rob.scala:339:30
  wire        T_28311_R6_data;	// rob.scala:339:30
  wire        T_28311_R7_data;	// rob.scala:339:30
  wire        T_28311_R8_data;	// rob.scala:339:30
  wire        T_28311_R9_data;	// rob.scala:339:30
  wire        T_28311_R10_data;	// rob.scala:339:30
  wire        T_28311_R11_data;	// rob.scala:339:30
  wire        T_28311_R12_data;	// rob.scala:339:30
  wire        T_28311_R13_data;	// rob.scala:339:30
  wire        T_28311_R14_data;	// rob.scala:339:30
  wire        T_28311_R15_data;	// rob.scala:339:30
  wire        T_28311_R16_data;	// rob.scala:339:30
  wire        T_28311_R17_data;	// rob.scala:339:30
  wire        T_28311_R18_data;	// rob.scala:339:30
  wire        T_28311_R19_data;	// rob.scala:339:30
  wire        T_28311_R20_data;	// rob.scala:339:30
  wire        T_28311_R21_data;	// rob.scala:339:30
  wire        T_28311_R22_data;	// rob.scala:339:30
  wire        T_28311_R23_data;	// rob.scala:339:30
  wire        T_28311_R24_data;	// rob.scala:339:30
  wire        T_23710_R0_data;	// rob.scala:335:30
  wire        T_23710_R1_data;	// rob.scala:335:30
  wire        T_23710_R2_data;	// rob.scala:335:30
  wire        T_23710_R3_data;	// rob.scala:335:30
  wire        T_23710_R4_data;	// rob.scala:335:30
  wire        T_23710_R5_data;	// rob.scala:335:30
  wire        T_23710_R6_data;	// rob.scala:335:30
  wire        T_23710_R7_data;	// rob.scala:335:30
  wire        T_23710_R8_data;	// rob.scala:335:30
  wire        T_23710_R9_data;	// rob.scala:335:30
  wire        T_23710_R10_data;	// rob.scala:335:30
  wire        T_23710_R11_data;	// rob.scala:335:30
  wire        T_23710_R12_data;	// rob.scala:335:30
  wire        T_23710_R13_data;	// rob.scala:335:30
  wire        T_23710_R14_data;	// rob.scala:335:30
  wire        T_23710_R15_data;	// rob.scala:335:30
  wire        T_23710_R16_data;	// rob.scala:335:30
  wire        T_23710_R17_data;	// rob.scala:335:30
  wire        T_23710_R18_data;	// rob.scala:335:30
  wire        T_23710_R19_data;	// rob.scala:335:30
  wire        T_23710_R20_data;	// rob.scala:335:30
  wire        T_23710_R21_data;	// rob.scala:335:30
  wire        T_23710_R22_data;	// rob.scala:335:30
  wire        T_23710_R23_data;	// rob.scala:335:30
  wire        T_23710_R24_data;	// rob.scala:335:30
  wire        row_metadata_has_brorjalr_R0_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R1_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R2_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R3_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R4_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R5_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R6_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R7_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R8_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R9_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R10_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R11_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R12_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R13_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R14_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R15_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R16_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R17_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R18_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R19_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R20_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R21_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R22_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R23_data;	// rob.scala:296:38
  wire        row_metadata_has_brorjalr_R24_data;	// rob.scala:296:38
  wire [4:0]  row_metadata_brob_idx_R2_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R3_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R4_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R5_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R6_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R7_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R8_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R9_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R10_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R11_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R12_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R13_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R14_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R15_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R16_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R17_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R18_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R19_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R20_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R21_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R22_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R23_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R24_data;	// rob.scala:295:35
  wire [4:0]  row_metadata_brob_idx_R25_data;	// rob.scala:295:35
  wire [36:0] T_23558_R0_data;	// rob.scala:894:22
  wire [36:0] T_23558_R1_data;	// rob.scala:894:22
  wire [36:0] T_23558_R2_data;	// rob.scala:894:22
  wire [36:0] T_23558_R3_data;	// rob.scala:894:22
  wire [36:0] T_23558_R4_data;	// rob.scala:894:22
  wire [36:0] T_23558_R5_data;	// rob.scala:894:22
  wire [36:0] T_23558_R6_data;	// rob.scala:894:22
  wire [36:0] T_23558_R7_data;	// rob.scala:894:22
  wire [36:0] T_23558_R8_data;	// rob.scala:894:22
  wire [36:0] T_23558_R9_data;	// rob.scala:894:22
  wire [36:0] T_23558_R10_data;	// rob.scala:894:22
  wire [36:0] T_23558_R11_data;	// rob.scala:894:22
  wire [36:0] T_23558_R12_data;	// rob.scala:894:22
  wire [36:0] T_23558_R13_data;	// rob.scala:894:22
  wire [36:0] T_23558_R14_data;	// rob.scala:894:22
  wire [36:0] T_23558_R15_data;	// rob.scala:894:22
  wire [36:0] T_23558_R16_data;	// rob.scala:894:22
  wire [36:0] T_23558_R17_data;	// rob.scala:894:22
  wire [36:0] T_23558_R18_data;	// rob.scala:894:22
  wire [36:0] T_23558_R19_data;	// rob.scala:894:22
  wire [36:0] T_23558_R20_data;	// rob.scala:894:22
  wire [36:0] T_23558_R21_data;	// rob.scala:894:22
  wire [36:0] T_23558_R22_data;	// rob.scala:894:22
  wire [36:0] T_23558_R23_data;	// rob.scala:894:22
  wire [36:0] T_23558_R24_data;	// rob.scala:894:22
  wire [36:0] T_23558_R25_data;	// rob.scala:894:22
  wire [36:0] T_23558_R26_data;	// rob.scala:894:22
  wire [36:0] T_23558_R27_data;	// rob.scala:894:22
  wire [36:0] T_23558_R28_data;	// rob.scala:894:22
  wire [36:0] T_23558_R29_data;	// rob.scala:894:22
  wire [36:0] T_23558_R30_data;	// rob.scala:894:22
  wire [36:0] T_23558_R31_data;	// rob.scala:894:22
  wire [36:0] T_23558_R32_data;	// rob.scala:894:22
  wire [36:0] T_23558_R33_data;	// rob.scala:894:22
  wire [36:0] T_23558_R34_data;	// rob.scala:894:22
  wire [36:0] T_23558_R35_data;	// rob.scala:894:22
  wire [36:0] T_23558_R36_data;	// rob.scala:894:22
  wire [36:0] T_23558_R37_data;	// rob.scala:894:22
  wire [36:0] T_23558_R38_data;	// rob.scala:894:22
  wire [36:0] T_23558_R39_data;	// rob.scala:894:22
  wire [36:0] T_23558_R40_data;	// rob.scala:894:22
  wire [36:0] T_23558_R41_data;	// rob.scala:894:22
  wire [36:0] T_23558_R42_data;	// rob.scala:894:22
  wire [36:0] T_23558_R43_data;	// rob.scala:894:22
  wire [36:0] T_23558_R44_data;	// rob.scala:894:22
  wire [36:0] T_23558_R45_data;	// rob.scala:894:22
  wire [36:0] T_23558_R46_data;	// rob.scala:894:22
  wire [36:0] T_23558_R47_data;	// rob.scala:894:22
  wire [36:0] T_23558_R48_data;	// rob.scala:894:22
  wire [36:0] T_23558_R49_data;	// rob.scala:894:22
  wire [36:0] T_23555_R0_data;	// rob.scala:893:22
  wire [36:0] T_23555_R1_data;	// rob.scala:893:22
  wire [36:0] T_23555_R2_data;	// rob.scala:893:22
  wire [36:0] T_23555_R3_data;	// rob.scala:893:22
  wire [36:0] T_23555_R4_data;	// rob.scala:893:22
  wire [36:0] T_23555_R5_data;	// rob.scala:893:22
  wire [36:0] T_23555_R6_data;	// rob.scala:893:22
  wire [36:0] T_23555_R7_data;	// rob.scala:893:22
  wire [36:0] T_23555_R8_data;	// rob.scala:893:22
  wire [36:0] T_23555_R9_data;	// rob.scala:893:22
  wire [36:0] T_23555_R10_data;	// rob.scala:893:22
  wire [36:0] T_23555_R11_data;	// rob.scala:893:22
  wire [36:0] T_23555_R12_data;	// rob.scala:893:22
  wire [36:0] T_23555_R13_data;	// rob.scala:893:22
  wire [36:0] T_23555_R14_data;	// rob.scala:893:22
  wire [36:0] T_23555_R15_data;	// rob.scala:893:22
  wire [36:0] T_23555_R16_data;	// rob.scala:893:22
  wire [36:0] T_23555_R17_data;	// rob.scala:893:22
  wire [36:0] T_23555_R18_data;	// rob.scala:893:22
  wire [36:0] T_23555_R19_data;	// rob.scala:893:22
  wire [36:0] T_23555_R20_data;	// rob.scala:893:22
  wire [36:0] T_23555_R21_data;	// rob.scala:893:22
  wire [36:0] T_23555_R22_data;	// rob.scala:893:22
  wire [36:0] T_23555_R23_data;	// rob.scala:893:22
  wire [36:0] T_23555_R24_data;	// rob.scala:893:22
  wire [36:0] T_23555_R25_data;	// rob.scala:893:22
  wire [36:0] T_23555_R26_data;	// rob.scala:893:22
  wire [36:0] T_23555_R27_data;	// rob.scala:893:22
  wire [36:0] T_23555_R28_data;	// rob.scala:893:22
  wire [36:0] T_23555_R29_data;	// rob.scala:893:22
  wire [36:0] T_23555_R30_data;	// rob.scala:893:22
  wire [36:0] T_23555_R31_data;	// rob.scala:893:22
  wire [36:0] T_23555_R32_data;	// rob.scala:893:22
  wire [36:0] T_23555_R33_data;	// rob.scala:893:22
  wire [36:0] T_23555_R34_data;	// rob.scala:893:22
  wire [36:0] T_23555_R35_data;	// rob.scala:893:22
  wire [36:0] T_23555_R36_data;	// rob.scala:893:22
  wire [36:0] T_23555_R37_data;	// rob.scala:893:22
  wire [36:0] T_23555_R38_data;	// rob.scala:893:22
  wire [36:0] T_23555_R39_data;	// rob.scala:893:22
  wire [36:0] T_23555_R40_data;	// rob.scala:893:22
  wire [36:0] T_23555_R41_data;	// rob.scala:893:22
  wire [36:0] T_23555_R42_data;	// rob.scala:893:22
  wire [36:0] T_23555_R43_data;	// rob.scala:893:22
  wire [36:0] T_23555_R44_data;	// rob.scala:893:22
  wire [36:0] T_23555_R45_data;	// rob.scala:893:22
  wire [36:0] T_23555_R46_data;	// rob.scala:893:22
  wire [36:0] T_23555_R47_data;	// rob.scala:893:22
  wire [36:0] T_23555_R48_data;	// rob.scala:893:22
  wire [36:0] T_23555_R49_data;	// rob.scala:893:22
  reg         casez_tmp;	// rob.scala:355:47
  reg         casez_tmp_2;	// rob.scala:433:51
  reg         casez_tmp_3;	// rob.scala:451:58
  reg         casez_tmp_4;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_5;	// rob.scala:453:59
  reg  [8:0]  casez_tmp_6;	// rob.scala:453:59
  reg  [31:0] casez_tmp_7;	// rob.scala:453:59
  reg  [39:0] casez_tmp_8;	// rob.scala:453:59
  reg  [7:0]  casez_tmp_9;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_10;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_11;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_12;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_13;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_14;	// rob.scala:453:59
  reg         casez_tmp_15;	// rob.scala:453:59
  reg         casez_tmp_16;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_17;	// rob.scala:453:59
  reg         casez_tmp_18;	// rob.scala:453:59
  reg         casez_tmp_19;	// rob.scala:453:59
  reg         casez_tmp_20;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_21;	// rob.scala:453:59
  reg         casez_tmp_22;	// rob.scala:453:59
  reg         casez_tmp_23;	// rob.scala:453:59
  reg         casez_tmp_24;	// rob.scala:453:59
  reg         casez_tmp_25;	// rob.scala:453:59
  reg         casez_tmp_26;	// rob.scala:453:59
  reg         casez_tmp_27;	// rob.scala:453:59
  reg  [7:0]  casez_tmp_28;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_29;	// rob.scala:453:59
  reg         casez_tmp_30;	// rob.scala:453:59
  reg         casez_tmp_31;	// rob.scala:453:59
  reg         casez_tmp_32;	// rob.scala:453:59
  reg         casez_tmp_33;	// rob.scala:453:59
  reg         casez_tmp_34;	// rob.scala:453:59
  reg         casez_tmp_35;	// rob.scala:453:59
  reg         casez_tmp_36;	// rob.scala:453:59
  reg         casez_tmp_37;	// rob.scala:453:59
  reg         casez_tmp_38;	// rob.scala:453:59
  reg         casez_tmp_39;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_40;	// rob.scala:453:59
  reg  [19:0] casez_tmp_41;	// rob.scala:453:59
  reg  [11:0] casez_tmp_42;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_43;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_44;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_45;	// rob.scala:453:59
  reg  [4:0]  casez_tmp_46;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_47;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_48;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_49;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_50;	// rob.scala:453:59
  reg         casez_tmp_51;	// rob.scala:453:59
  reg         casez_tmp_52;	// rob.scala:453:59
  reg         casez_tmp_53;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_54;	// rob.scala:453:59
  reg         casez_tmp_55;	// rob.scala:453:59
  reg  [63:0] casez_tmp_56;	// rob.scala:453:59
  reg         casez_tmp_57;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_58;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_59;	// rob.scala:453:59
  reg         casez_tmp_60;	// rob.scala:453:59
  reg         casez_tmp_61;	// rob.scala:453:59
  reg         casez_tmp_62;	// rob.scala:453:59
  reg         casez_tmp_63;	// rob.scala:453:59
  reg         casez_tmp_64;	// rob.scala:453:59
  reg         casez_tmp_65;	// rob.scala:453:59
  reg         casez_tmp_66;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_67;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_68;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_69;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_70;	// rob.scala:453:59
  reg         casez_tmp_71;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_72;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_73;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_74;	// rob.scala:453:59
  reg         casez_tmp_75;	// rob.scala:453:59
  reg         casez_tmp_76;	// rob.scala:453:59
  reg         casez_tmp_77;	// rob.scala:453:59
  reg         casez_tmp_78;	// rob.scala:453:59
  reg         casez_tmp_79;	// rob.scala:453:59
  reg  [31:0] casez_tmp_80;	// rob.scala:453:59
  reg         casez_tmp_81;	// rob.scala:507:28
  reg         casez_tmp_82;	// rob.scala:507:28
  reg  [63:0] casez_tmp_83;	// rob.scala:507:28
  reg         casez_tmp_84;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_85;	// rob.scala:538:75
  reg         casez_tmp_86;	// rob.scala:538:75
  reg         casez_tmp_87;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_88;	// rob.scala:538:75
  reg         casez_tmp_89;	// rob.scala:538:75
  reg         casez_tmp_90;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_91;	// rob.scala:538:75
  reg         casez_tmp_92;	// rob.scala:538:75
  reg         casez_tmp_93;	// rob.scala:355:47
  reg         casez_tmp_94;	// rob.scala:433:51
  reg         casez_tmp_95;	// rob.scala:451:58
  reg         casez_tmp_96;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_97;	// rob.scala:453:59
  reg  [8:0]  casez_tmp_98;	// rob.scala:453:59
  reg  [31:0] casez_tmp_99;	// rob.scala:453:59
  reg  [39:0] casez_tmp_100;	// rob.scala:453:59
  reg  [7:0]  casez_tmp_101;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_102;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_103;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_104;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_105;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_106;	// rob.scala:453:59
  reg         casez_tmp_107;	// rob.scala:453:59
  reg         casez_tmp_108;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_109;	// rob.scala:453:59
  reg         casez_tmp_110;	// rob.scala:453:59
  reg         casez_tmp_111;	// rob.scala:453:59
  reg         casez_tmp_112;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_113;	// rob.scala:453:59
  reg         casez_tmp_114;	// rob.scala:453:59
  reg         casez_tmp_115;	// rob.scala:453:59
  reg         casez_tmp_116;	// rob.scala:453:59
  reg         casez_tmp_117;	// rob.scala:453:59
  reg         casez_tmp_118;	// rob.scala:453:59
  reg         casez_tmp_119;	// rob.scala:453:59
  reg  [7:0]  casez_tmp_120;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_121;	// rob.scala:453:59
  reg         casez_tmp_122;	// rob.scala:453:59
  reg         casez_tmp_123;	// rob.scala:453:59
  reg         casez_tmp_124;	// rob.scala:453:59
  reg         casez_tmp_125;	// rob.scala:453:59
  reg         casez_tmp_126;	// rob.scala:453:59
  reg         casez_tmp_127;	// rob.scala:453:59
  reg         casez_tmp_128;	// rob.scala:453:59
  reg         casez_tmp_129;	// rob.scala:453:59
  reg         casez_tmp_130;	// rob.scala:453:59
  reg         casez_tmp_131;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_132;	// rob.scala:453:59
  reg  [19:0] casez_tmp_133;	// rob.scala:453:59
  reg  [11:0] casez_tmp_134;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_135;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_136;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_137;	// rob.scala:453:59
  reg  [4:0]  casez_tmp_138;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_139;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_140;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_141;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_142;	// rob.scala:453:59
  reg         casez_tmp_143;	// rob.scala:453:59
  reg         casez_tmp_144;	// rob.scala:453:59
  reg         casez_tmp_145;	// rob.scala:453:59
  reg  [6:0]  casez_tmp_146;	// rob.scala:453:59
  reg         casez_tmp_147;	// rob.scala:453:59
  reg  [63:0] casez_tmp_148;	// rob.scala:453:59
  reg         casez_tmp_149;	// rob.scala:453:59
  reg  [3:0]  casez_tmp_150;	// rob.scala:453:59
  reg  [2:0]  casez_tmp_151;	// rob.scala:453:59
  reg         casez_tmp_152;	// rob.scala:453:59
  reg         casez_tmp_153;	// rob.scala:453:59
  reg         casez_tmp_154;	// rob.scala:453:59
  reg         casez_tmp_155;	// rob.scala:453:59
  reg         casez_tmp_156;	// rob.scala:453:59
  reg         casez_tmp_157;	// rob.scala:453:59
  reg         casez_tmp_158;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_159;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_160;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_161;	// rob.scala:453:59
  reg  [5:0]  casez_tmp_162;	// rob.scala:453:59
  reg         casez_tmp_163;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_164;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_165;	// rob.scala:453:59
  reg  [1:0]  casez_tmp_166;	// rob.scala:453:59
  reg         casez_tmp_167;	// rob.scala:453:59
  reg         casez_tmp_168;	// rob.scala:453:59
  reg         casez_tmp_169;	// rob.scala:453:59
  reg         casez_tmp_170;	// rob.scala:453:59
  reg         casez_tmp_171;	// rob.scala:453:59
  reg  [31:0] casez_tmp_172;	// rob.scala:453:59
  reg         casez_tmp_173;	// rob.scala:507:28
  reg         casez_tmp_174;	// rob.scala:507:28
  reg  [63:0] casez_tmp_175;	// rob.scala:507:28
  reg         casez_tmp_176;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_177;	// rob.scala:538:75
  reg         casez_tmp_178;	// rob.scala:538:75
  reg         casez_tmp_179;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_180;	// rob.scala:538:75
  reg         casez_tmp_181;	// rob.scala:538:75
  reg         casez_tmp_182;	// rob.scala:536:22
  reg  [6:0]  casez_tmp_183;	// rob.scala:538:75
  reg         casez_tmp_184;	// rob.scala:538:75
  reg  [7:0]  casez_tmp_185;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_186;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_187;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_188;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_189;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_190;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_191;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_192;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_193;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_194;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_195;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_196;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_197;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_198;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_199;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_200;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_201;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_202;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_203;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_204;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_205;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_206;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_207;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_208;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_209;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_210;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_211;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_212;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_213;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_214;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_215;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_216;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_217;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_218;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_219;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_220;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_221;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_222;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_223;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_224;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_225;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_226;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_227;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_228;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_229;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_230;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_231;	// rob.scala:1048:21
  reg  [7:0]  casez_tmp_232;	// rob.scala:1048:21
  reg  [1:0]  rob_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
  reg  [4:0]  rob_head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:5
  reg  [4:0]  rob_tail;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:14:5
  reg         r_xcpt_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:36:5
  reg         r_xcpt_uop_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [8:0]  r_xcpt_uop_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [31:0] r_xcpt_uop_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [39:0] r_xcpt_uop_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [7:0]  r_xcpt_uop_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [3:0]  r_xcpt_uop_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [3:0]  r_xcpt_uop_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [7:0]  r_xcpt_uop_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [19:0] r_xcpt_uop_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [11:0] r_xcpt_uop_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [5:0]  r_xcpt_uop_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [3:0]  r_xcpt_uop_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [3:0]  r_xcpt_uop_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [4:0]  r_xcpt_uop_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [6:0]  r_xcpt_uop_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [6:0]  r_xcpt_uop_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [6:0]  r_xcpt_uop_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [6:0]  r_xcpt_uop_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [6:0]  r_xcpt_uop_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [63:0] r_xcpt_uop_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [3:0]  r_xcpt_uop_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [2:0]  r_xcpt_uop_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [5:0]  r_xcpt_uop_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [5:0]  r_xcpt_uop_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [5:0]  r_xcpt_uop_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [5:0]  r_xcpt_uop_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [1:0]  r_xcpt_uop_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg         r_xcpt_uop_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [63:0] r_xcpt_uop_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [31:0] r_xcpt_uop_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
  reg  [39:0] r_xcpt_badvaddr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:38:5
  reg         r_partial_row;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:125:5
  reg         T_23706_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_8;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_9;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_10;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_11;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_12;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_13;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_14;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_15;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_16;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_17;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_18;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_19;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_20;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_21;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_22;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_23706_23;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
  reg         T_26182_0_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_0_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_0_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_0_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_0_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_0_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_0_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_0_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_0_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_0_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_0_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_0_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_0_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_0_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_0_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_0_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_0_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_0_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_0_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_0_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_0_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_0_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_0_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_0_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_0_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_0_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_0_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_0_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_0_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_0_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_1_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_1_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_1_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_1_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_1_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_1_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_1_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_1_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_1_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_1_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_1_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_1_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_1_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_1_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_1_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_1_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_1_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_1_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_1_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_1_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_1_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_1_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_1_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_1_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_1_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_1_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_1_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_1_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_1_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_2_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_2_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_2_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_2_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_2_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_2_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_2_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_2_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_2_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_2_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_2_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_2_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_2_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_2_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_2_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_2_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_2_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_2_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_2_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_2_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_2_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_2_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_2_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_2_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_2_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_2_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_2_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_2_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_2_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_3_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_3_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_3_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_3_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_3_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_3_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_3_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_3_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_3_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_3_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_3_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_3_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_3_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_3_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_3_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_3_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_3_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_3_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_3_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_3_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_3_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_3_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_3_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_3_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_3_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_3_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_3_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_3_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_3_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_4_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_4_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_4_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_4_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_4_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_4_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_4_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_4_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_4_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_4_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_4_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_4_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_4_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_4_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_4_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_4_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_4_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_4_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_4_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_4_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_4_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_4_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_4_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_4_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_4_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_4_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_4_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_4_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_4_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_5_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_5_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_5_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_5_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_5_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_5_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_5_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_5_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_5_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_5_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_5_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_5_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_5_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_5_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_5_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_5_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_5_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_5_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_5_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_5_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_5_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_5_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_5_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_5_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_5_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_5_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_5_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_5_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_5_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_6_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_6_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_6_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_6_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_6_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_6_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_6_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_6_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_6_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_6_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_6_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_6_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_6_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_6_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_6_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_6_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_6_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_6_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_6_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_6_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_6_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_6_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_6_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_6_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_6_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_6_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_6_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_6_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_6_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_7_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_7_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_7_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_7_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_7_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_7_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_7_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_7_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_7_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_7_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_7_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_7_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_7_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_7_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_7_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_7_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_7_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_7_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_7_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_7_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_7_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_7_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_7_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_7_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_7_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_7_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_7_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_7_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_7_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_8_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_8_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_8_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_8_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_8_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_8_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_8_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_8_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_8_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_8_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_8_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_8_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_8_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_8_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_8_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_8_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_8_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_8_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_8_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_8_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_8_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_8_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_8_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_8_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_8_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_8_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_8_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_8_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_8_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_9_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_9_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_9_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_9_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_9_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_9_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_9_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_9_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_9_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_9_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_9_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_9_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_9_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_9_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_9_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_9_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_9_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_9_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_9_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_9_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_9_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_9_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_9_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_9_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_9_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_9_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_9_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_9_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_9_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_10_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_10_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_10_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_10_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_10_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_10_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_10_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_10_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_10_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_10_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_10_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_10_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_10_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_10_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_10_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_10_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_10_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_10_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_10_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_10_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_10_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_10_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_10_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_10_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_10_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_10_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_10_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_10_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_10_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_11_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_11_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_11_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_11_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_11_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_11_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_11_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_11_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_11_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_11_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_11_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_11_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_11_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_11_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_11_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_11_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_11_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_11_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_11_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_11_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_11_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_11_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_11_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_11_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_11_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_11_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_11_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_11_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_11_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_12_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_12_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_12_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_12_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_12_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_12_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_12_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_12_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_12_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_12_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_12_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_12_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_12_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_12_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_12_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_12_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_12_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_12_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_12_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_12_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_12_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_12_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_12_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_12_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_12_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_12_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_12_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_12_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_12_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_13_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_13_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_13_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_13_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_13_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_13_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_13_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_13_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_13_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_13_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_13_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_13_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_13_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_13_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_13_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_13_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_13_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_13_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_13_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_13_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_13_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_13_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_13_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_13_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_13_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_13_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_13_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_13_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_13_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_14_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_14_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_14_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_14_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_14_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_14_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_14_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_14_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_14_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_14_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_14_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_14_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_14_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_14_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_14_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_14_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_14_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_14_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_14_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_14_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_14_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_14_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_14_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_14_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_14_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_14_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_14_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_14_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_14_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_15_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_15_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_15_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_15_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_15_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_15_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_15_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_15_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_15_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_15_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_15_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_15_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_15_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_15_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_15_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_15_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_15_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_15_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_15_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_15_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_15_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_15_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_15_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_15_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_15_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_15_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_15_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_15_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_15_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_16_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_16_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_16_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_16_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_16_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_16_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_16_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_16_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_16_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_16_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_16_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_16_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_16_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_16_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_16_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_16_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_16_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_16_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_16_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_16_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_16_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_16_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_16_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_16_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_16_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_16_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_16_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_16_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_16_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_17_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_17_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_17_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_17_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_17_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_17_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_17_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_17_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_17_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_17_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_17_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_17_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_17_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_17_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_17_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_17_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_17_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_17_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_17_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_17_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_17_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_17_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_17_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_17_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_17_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_17_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_17_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_17_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_17_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_18_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_18_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_18_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_18_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_18_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_18_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_18_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_18_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_18_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_18_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_18_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_18_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_18_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_18_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_18_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_18_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_18_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_18_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_18_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_18_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_18_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_18_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_18_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_18_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_18_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_18_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_18_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_18_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_18_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_19_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_19_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_19_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_19_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_19_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_19_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_19_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_19_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_19_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_19_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_19_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_19_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_19_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_19_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_19_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_19_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_19_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_19_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_19_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_19_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_19_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_19_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_19_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_19_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_19_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_19_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_19_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_19_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_19_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_20_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_20_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_20_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_20_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_20_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_20_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_20_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_20_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_20_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_20_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_20_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_20_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_20_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_20_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_20_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_20_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_20_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_20_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_20_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_20_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_20_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_20_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_20_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_20_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_20_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_20_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_20_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_20_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_20_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_21_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_21_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_21_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_21_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_21_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_21_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_21_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_21_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_21_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_21_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_21_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_21_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_21_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_21_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_21_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_21_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_21_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_21_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_21_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_21_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_21_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_21_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_21_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_21_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_21_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_21_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_21_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_21_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_21_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_22_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_22_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_22_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_22_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_22_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_22_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_22_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_22_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_22_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_22_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_22_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_22_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_22_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_22_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_22_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_22_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_22_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_22_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_22_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_22_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_22_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_22_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_22_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_22_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_22_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_22_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_22_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_22_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_22_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [8:0]  T_26182_23_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_23_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [39:0] T_26182_23_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_23_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_23_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_23_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [7:0]  T_26182_23_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [19:0] T_26182_23_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [11:0] T_26182_23_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_23_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_23_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_23_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [4:0]  T_26182_23_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_23_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_23_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_23_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_23_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [6:0]  T_26182_23_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_23_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [3:0]  T_26182_23_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [2:0]  T_26182_23_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_23_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_23_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_23_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [5:0]  T_26182_23_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [1:0]  T_26182_23_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_26182_23_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [63:0] T_26182_23_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg  [31:0] T_26182_23_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
  reg         T_35634_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_8;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_9;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_10;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_11;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_12;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_13;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_14;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_15;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_16;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_17;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_18;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_19;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_20;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_21;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_22;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_35634_23;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
  reg         T_38110_0_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_0_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_0_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_0_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_0_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_0_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_0_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_0_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_0_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_0_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_0_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_0_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_0_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_0_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_0_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_0_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_0_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_0_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_0_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_0_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_0_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_0_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_0_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_0_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_0_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_0_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_0_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_0_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_0_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_0_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_1_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_1_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_1_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_1_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_1_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_1_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_1_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_1_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_1_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_1_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_1_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_1_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_1_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_1_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_1_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_1_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_1_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_1_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_1_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_1_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_1_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_1_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_1_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_1_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_1_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_1_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_1_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_1_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_1_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_2_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_2_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_2_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_2_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_2_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_2_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_2_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_2_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_2_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_2_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_2_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_2_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_2_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_2_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_2_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_2_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_2_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_2_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_2_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_2_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_2_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_2_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_2_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_2_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_2_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_2_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_2_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_2_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_2_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_3_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_3_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_3_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_3_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_3_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_3_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_3_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_3_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_3_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_3_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_3_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_3_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_3_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_3_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_3_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_3_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_3_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_3_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_3_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_3_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_3_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_3_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_3_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_3_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_3_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_3_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_3_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_3_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_3_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_4_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_4_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_4_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_4_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_4_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_4_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_4_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_4_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_4_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_4_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_4_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_4_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_4_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_4_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_4_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_4_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_4_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_4_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_4_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_4_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_4_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_4_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_4_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_4_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_4_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_4_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_4_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_4_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_4_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_5_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_5_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_5_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_5_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_5_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_5_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_5_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_5_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_5_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_5_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_5_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_5_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_5_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_5_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_5_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_5_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_5_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_5_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_5_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_5_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_5_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_5_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_5_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_5_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_5_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_5_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_5_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_5_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_5_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_6_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_6_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_6_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_6_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_6_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_6_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_6_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_6_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_6_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_6_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_6_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_6_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_6_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_6_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_6_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_6_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_6_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_6_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_6_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_6_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_6_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_6_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_6_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_6_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_6_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_6_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_6_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_6_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_6_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_7_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_7_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_7_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_7_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_7_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_7_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_7_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_7_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_7_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_7_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_7_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_7_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_7_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_7_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_7_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_7_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_7_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_7_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_7_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_7_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_7_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_7_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_7_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_7_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_7_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_7_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_7_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_7_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_7_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_8_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_8_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_8_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_8_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_8_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_8_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_8_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_8_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_8_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_8_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_8_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_8_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_8_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_8_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_8_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_8_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_8_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_8_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_8_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_8_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_8_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_8_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_8_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_8_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_8_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_8_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_8_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_8_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_8_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_9_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_9_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_9_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_9_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_9_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_9_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_9_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_9_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_9_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_9_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_9_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_9_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_9_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_9_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_9_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_9_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_9_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_9_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_9_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_9_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_9_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_9_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_9_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_9_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_9_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_9_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_9_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_9_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_9_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_10_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_10_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_10_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_10_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_10_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_10_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_10_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_10_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_10_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_10_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_10_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_10_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_10_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_10_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_10_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_10_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_10_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_10_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_10_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_10_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_10_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_10_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_10_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_10_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_10_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_10_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_10_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_10_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_10_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_11_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_11_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_11_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_11_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_11_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_11_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_11_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_11_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_11_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_11_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_11_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_11_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_11_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_11_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_11_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_11_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_11_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_11_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_11_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_11_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_11_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_11_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_11_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_11_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_11_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_11_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_11_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_11_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_11_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_12_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_12_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_12_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_12_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_12_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_12_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_12_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_12_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_12_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_12_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_12_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_12_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_12_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_12_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_12_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_12_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_12_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_12_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_12_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_12_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_12_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_12_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_12_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_12_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_12_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_12_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_12_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_12_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_12_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_13_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_13_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_13_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_13_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_13_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_13_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_13_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_13_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_13_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_13_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_13_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_13_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_13_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_13_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_13_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_13_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_13_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_13_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_13_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_13_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_13_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_13_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_13_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_13_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_13_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_13_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_13_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_13_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_13_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_14_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_14_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_14_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_14_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_14_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_14_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_14_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_14_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_14_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_14_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_14_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_14_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_14_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_14_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_14_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_14_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_14_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_14_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_14_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_14_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_14_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_14_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_14_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_14_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_14_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_14_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_14_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_14_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_14_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_15_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_15_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_15_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_15_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_15_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_15_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_15_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_15_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_15_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_15_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_15_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_15_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_15_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_15_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_15_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_15_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_15_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_15_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_15_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_15_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_15_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_15_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_15_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_15_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_15_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_15_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_15_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_15_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_15_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_16_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_16_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_16_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_16_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_16_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_16_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_16_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_16_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_16_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_16_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_16_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_16_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_16_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_16_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_16_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_16_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_16_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_16_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_16_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_16_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_16_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_16_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_16_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_16_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_16_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_16_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_16_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_16_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_16_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_17_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_17_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_17_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_17_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_17_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_17_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_17_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_17_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_17_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_17_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_17_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_17_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_17_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_17_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_17_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_17_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_17_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_17_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_17_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_17_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_17_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_17_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_17_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_17_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_17_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_17_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_17_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_17_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_17_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_18_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_18_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_18_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_18_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_18_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_18_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_18_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_18_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_18_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_18_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_18_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_18_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_18_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_18_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_18_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_18_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_18_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_18_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_18_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_18_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_18_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_18_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_18_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_18_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_18_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_18_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_18_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_18_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_18_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_19_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_19_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_19_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_19_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_19_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_19_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_19_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_19_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_19_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_19_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_19_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_19_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_19_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_19_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_19_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_19_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_19_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_19_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_19_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_19_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_19_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_19_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_19_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_19_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_19_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_19_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_19_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_19_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_19_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_20_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_20_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_20_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_20_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_20_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_20_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_20_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_20_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_20_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_20_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_20_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_20_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_20_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_20_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_20_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_20_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_20_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_20_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_20_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_20_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_20_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_20_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_20_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_20_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_20_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_20_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_20_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_20_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_20_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_21_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_21_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_21_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_21_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_21_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_21_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_21_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_21_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_21_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_21_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_21_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_21_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_21_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_21_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_21_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_21_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_21_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_21_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_21_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_21_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_21_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_21_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_21_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_21_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_21_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_21_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_21_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_21_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_21_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_22_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_22_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_22_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_22_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_22_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_22_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_22_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_22_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_22_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_22_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_22_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_22_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_22_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_22_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_22_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_22_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_22_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_22_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_22_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_22_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_22_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_22_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_22_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_22_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_22_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_22_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_22_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_22_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_22_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [8:0]  T_38110_23_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_23_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [39:0] T_38110_23_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_23_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_23_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_23_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [7:0]  T_38110_23_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [19:0] T_38110_23_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [11:0] T_38110_23_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_23_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_23_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_23_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [4:0]  T_38110_23_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_23_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_23_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_23_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_23_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [6:0]  T_38110_23_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_23_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [3:0]  T_38110_23_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [2:0]  T_38110_23_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_23_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_23_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_23_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [5:0]  T_38110_23_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [1:0]  T_38110_23_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_38110_23_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [63:0] T_38110_23_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg  [31:0] T_38110_23_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
  reg         T_47576;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2940:5
  reg         T_47616;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2978:5

  wire _T_23559 = io_dis_valids_0 | io_dis_valids_1;	// rob.scala:260:32
  wire [36:0] _io_dis_uops_0_pc_39to3 = io_dis_uops_0_pc[39:3];	// rob.scala:931:42
  wire _T_23563 = rob_tail[0];	// rob.scala:192:32, :932:25
  wire [3:0] _rob_tail_4to1 = rob_tail[4:1];	// rob.scala:192:32, :934:29
  wire [4:0] _io_get_pc_rob_idx_5to1 = io_get_pc_rob_idx[5:1];	// rob.scala:222:27
  wire _io_get_pc_rob_idx_1 = io_get_pc_rob_idx[1];	// rob.scala:913:37
  wire [3:0] _io_get_pc_rob_idx_5to2 = io_get_pc_rob_idx[5:2];	// rob.scala:913:58
  wire _rob_pc_hob_next_val = _T_1 | _T_0;	// rob.scala:273:51, :509:28
  wire _T_23652 = _T_23559 & io_dis_new_packet;	// rob.scala:297:36
  wire _T_23670 = io_dis_valids_0 & io_dis_uops_0_is_unique;	// rob.scala:322:24
  wire _T_23671 = io_dis_valids_1 & io_dis_uops_1_is_unique;	// rob.scala:322:24
  wire _T_23672 = _T_23670 | _T_23671;	// rob.scala:322:61
  always @(*) begin	// rob.scala:347:34, :355:47
    casez (rob_tail)	// rob.scala:192:32, :347:34, :355:47
      5'b00000:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b00001:
        casez_tmp = T_23706_1;	// rob.scala:347:34, :355:47
      5'b00010:
        casez_tmp = T_23706_2;	// rob.scala:347:34, :355:47
      5'b00011:
        casez_tmp = T_23706_3;	// rob.scala:347:34, :355:47
      5'b00100:
        casez_tmp = T_23706_4;	// rob.scala:347:34, :355:47
      5'b00101:
        casez_tmp = T_23706_5;	// rob.scala:347:34, :355:47
      5'b00110:
        casez_tmp = T_23706_6;	// rob.scala:347:34, :355:47
      5'b00111:
        casez_tmp = T_23706_7;	// rob.scala:347:34, :355:47
      5'b01000:
        casez_tmp = T_23706_8;	// rob.scala:347:34, :355:47
      5'b01001:
        casez_tmp = T_23706_9;	// rob.scala:347:34, :355:47
      5'b01010:
        casez_tmp = T_23706_10;	// rob.scala:347:34, :355:47
      5'b01011:
        casez_tmp = T_23706_11;	// rob.scala:347:34, :355:47
      5'b01100:
        casez_tmp = T_23706_12;	// rob.scala:347:34, :355:47
      5'b01101:
        casez_tmp = T_23706_13;	// rob.scala:347:34, :355:47
      5'b01110:
        casez_tmp = T_23706_14;	// rob.scala:347:34, :355:47
      5'b01111:
        casez_tmp = T_23706_15;	// rob.scala:347:34, :355:47
      5'b10000:
        casez_tmp = T_23706_16;	// rob.scala:347:34, :355:47
      5'b10001:
        casez_tmp = T_23706_17;	// rob.scala:347:34, :355:47
      5'b10010:
        casez_tmp = T_23706_18;	// rob.scala:347:34, :355:47
      5'b10011:
        casez_tmp = T_23706_19;	// rob.scala:347:34, :355:47
      5'b10100:
        casez_tmp = T_23706_20;	// rob.scala:347:34, :355:47
      5'b10101:
        casez_tmp = T_23706_21;	// rob.scala:347:34, :355:47
      5'b10110:
        casez_tmp = T_23706_22;	// rob.scala:347:34, :355:47
      5'b10111:
        casez_tmp = T_23706_23;	// rob.scala:347:34, :355:47
      5'b11000:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11001:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11010:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11011:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11100:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11101:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      5'b11110:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
      default:
        casez_tmp = T_23706_0;	// rob.scala:347:34, :355:47
    endcase	// rob.scala:192:32, :347:34, :355:47
  end // always @(*)
  wire [4:0] _io_wb_resps_0_bits_uop_rob_idx_5to1 = io_wb_resps_0_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_28590 = io_wb_resps_0_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_wb_resps_1_bits_uop_rob_idx_5to1 = io_wb_resps_1_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_28598 = io_wb_resps_1_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_wb_resps_2_bits_uop_rob_idx_5to1 = io_wb_resps_2_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_28606 = io_wb_resps_2_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire _T_28612 = io_lsu_clr_bsy_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_lsu_clr_bsy_rob_idx_5to1 = io_lsu_clr_bsy_rob_idx[5:1];	// rob.scala:222:27
  wire _T_29059 = io_fflags_0_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_fflags_0_bits_uop_rob_idx_5to1 = io_fflags_0_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_29066 = io_fflags_1_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_fflags_1_bits_uop_rob_idx_5to1 = io_fflags_1_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_29073 = io_lxcpt_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_lxcpt_bits_uop_rob_idx_5to1 = io_lxcpt_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  wire _T_29081 = io_bxcpt_bits_uop_rob_idx[0];	// rob.scala:227:38
  wire [4:0] _io_bxcpt_bits_uop_rob_idx_5to1 = io_bxcpt_bits_uop_rob_idx[5:1];	// rob.scala:222:27
  always @(*) begin	// rob.scala:433:51
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51
      5'b00000:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b00001:
        casez_tmp_2 = T_23706_1;	// rob.scala:347:34, :433:51
      5'b00010:
        casez_tmp_2 = T_23706_2;	// rob.scala:347:34, :433:51
      5'b00011:
        casez_tmp_2 = T_23706_3;	// rob.scala:347:34, :433:51
      5'b00100:
        casez_tmp_2 = T_23706_4;	// rob.scala:347:34, :433:51
      5'b00101:
        casez_tmp_2 = T_23706_5;	// rob.scala:347:34, :433:51
      5'b00110:
        casez_tmp_2 = T_23706_6;	// rob.scala:347:34, :433:51
      5'b00111:
        casez_tmp_2 = T_23706_7;	// rob.scala:347:34, :433:51
      5'b01000:
        casez_tmp_2 = T_23706_8;	// rob.scala:347:34, :433:51
      5'b01001:
        casez_tmp_2 = T_23706_9;	// rob.scala:347:34, :433:51
      5'b01010:
        casez_tmp_2 = T_23706_10;	// rob.scala:347:34, :433:51
      5'b01011:
        casez_tmp_2 = T_23706_11;	// rob.scala:347:34, :433:51
      5'b01100:
        casez_tmp_2 = T_23706_12;	// rob.scala:347:34, :433:51
      5'b01101:
        casez_tmp_2 = T_23706_13;	// rob.scala:347:34, :433:51
      5'b01110:
        casez_tmp_2 = T_23706_14;	// rob.scala:347:34, :433:51
      5'b01111:
        casez_tmp_2 = T_23706_15;	// rob.scala:347:34, :433:51
      5'b10000:
        casez_tmp_2 = T_23706_16;	// rob.scala:347:34, :433:51
      5'b10001:
        casez_tmp_2 = T_23706_17;	// rob.scala:347:34, :433:51
      5'b10010:
        casez_tmp_2 = T_23706_18;	// rob.scala:347:34, :433:51
      5'b10011:
        casez_tmp_2 = T_23706_19;	// rob.scala:347:34, :433:51
      5'b10100:
        casez_tmp_2 = T_23706_20;	// rob.scala:347:34, :433:51
      5'b10101:
        casez_tmp_2 = T_23706_21;	// rob.scala:347:34, :433:51
      5'b10110:
        casez_tmp_2 = T_23706_22;	// rob.scala:347:34, :433:51
      5'b10111:
        casez_tmp_2 = T_23706_23;	// rob.scala:347:34, :433:51
      5'b11000:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11001:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11010:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11011:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11100:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11101:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      5'b11110:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
      default:
        casez_tmp_2 = T_23706_0;	// rob.scala:347:34, :433:51
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51
  end // always @(*)
  wire _T_29090 = casez_tmp_2 & T_28311_R0_data;	// rob.scala:339:30, :433:51
  wire _T_29094 = casez_tmp_2 & ~T_23710_R0_data;	// rob.scala:335:30, :433:51, :439:{42,45}
  wire _T_29097 = rob_state == 2'h2;	// rob.scala:443:23
  wire [4:0] _T_2 = _T_29097 ? rob_tail : rob_head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :445:18
  always @(*) begin	// rob.scala:451:58
    casez (_T_2)	// rob.scala:451:58
      5'b00000:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b00001:
        casez_tmp_3 = T_23706_1;	// rob.scala:347:34, :451:58
      5'b00010:
        casez_tmp_3 = T_23706_2;	// rob.scala:347:34, :451:58
      5'b00011:
        casez_tmp_3 = T_23706_3;	// rob.scala:347:34, :451:58
      5'b00100:
        casez_tmp_3 = T_23706_4;	// rob.scala:347:34, :451:58
      5'b00101:
        casez_tmp_3 = T_23706_5;	// rob.scala:347:34, :451:58
      5'b00110:
        casez_tmp_3 = T_23706_6;	// rob.scala:347:34, :451:58
      5'b00111:
        casez_tmp_3 = T_23706_7;	// rob.scala:347:34, :451:58
      5'b01000:
        casez_tmp_3 = T_23706_8;	// rob.scala:347:34, :451:58
      5'b01001:
        casez_tmp_3 = T_23706_9;	// rob.scala:347:34, :451:58
      5'b01010:
        casez_tmp_3 = T_23706_10;	// rob.scala:347:34, :451:58
      5'b01011:
        casez_tmp_3 = T_23706_11;	// rob.scala:347:34, :451:58
      5'b01100:
        casez_tmp_3 = T_23706_12;	// rob.scala:347:34, :451:58
      5'b01101:
        casez_tmp_3 = T_23706_13;	// rob.scala:347:34, :451:58
      5'b01110:
        casez_tmp_3 = T_23706_14;	// rob.scala:347:34, :451:58
      5'b01111:
        casez_tmp_3 = T_23706_15;	// rob.scala:347:34, :451:58
      5'b10000:
        casez_tmp_3 = T_23706_16;	// rob.scala:347:34, :451:58
      5'b10001:
        casez_tmp_3 = T_23706_17;	// rob.scala:347:34, :451:58
      5'b10010:
        casez_tmp_3 = T_23706_18;	// rob.scala:347:34, :451:58
      5'b10011:
        casez_tmp_3 = T_23706_19;	// rob.scala:347:34, :451:58
      5'b10100:
        casez_tmp_3 = T_23706_20;	// rob.scala:347:34, :451:58
      5'b10101:
        casez_tmp_3 = T_23706_21;	// rob.scala:347:34, :451:58
      5'b10110:
        casez_tmp_3 = T_23706_22;	// rob.scala:347:34, :451:58
      5'b10111:
        casez_tmp_3 = T_23706_23;	// rob.scala:347:34, :451:58
      5'b11000:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11001:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11010:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11011:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11100:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11101:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      5'b11110:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
      default:
        casez_tmp_3 = T_23706_0;	// rob.scala:347:34, :451:58
    endcase	// rob.scala:451:58
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_4 = T_26182_1_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_4 = T_26182_2_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_4 = T_26182_3_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_4 = T_26182_4_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_4 = T_26182_5_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_4 = T_26182_6_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_4 = T_26182_7_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_4 = T_26182_8_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_4 = T_26182_9_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_4 = T_26182_10_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_4 = T_26182_11_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_4 = T_26182_12_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_4 = T_26182_13_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_4 = T_26182_14_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_4 = T_26182_15_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_4 = T_26182_16_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_4 = T_26182_17_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_4 = T_26182_18_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_4 = T_26182_19_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_4 = T_26182_20_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_4 = T_26182_21_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_4 = T_26182_22_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_4 = T_26182_23_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_4 = T_26182_0_valid;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_5 = T_26182_1_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_5 = T_26182_2_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_5 = T_26182_3_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_5 = T_26182_4_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_5 = T_26182_5_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_5 = T_26182_6_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_5 = T_26182_7_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_5 = T_26182_8_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_5 = T_26182_9_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_5 = T_26182_10_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_5 = T_26182_11_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_5 = T_26182_12_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_5 = T_26182_13_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_5 = T_26182_14_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_5 = T_26182_15_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_5 = T_26182_16_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_5 = T_26182_17_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_5 = T_26182_18_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_5 = T_26182_19_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_5 = T_26182_20_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_5 = T_26182_21_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_5 = T_26182_22_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_5 = T_26182_23_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_5 = T_26182_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_6 = T_26182_1_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_6 = T_26182_2_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_6 = T_26182_3_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_6 = T_26182_4_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_6 = T_26182_5_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_6 = T_26182_6_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_6 = T_26182_7_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_6 = T_26182_8_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_6 = T_26182_9_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_6 = T_26182_10_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_6 = T_26182_11_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_6 = T_26182_12_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_6 = T_26182_13_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_6 = T_26182_14_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_6 = T_26182_15_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_6 = T_26182_16_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_6 = T_26182_17_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_6 = T_26182_18_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_6 = T_26182_19_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_6 = T_26182_20_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_6 = T_26182_21_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_6 = T_26182_22_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_6 = T_26182_23_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_6 = T_26182_0_uopc;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_7 = T_26182_1_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_7 = T_26182_2_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_7 = T_26182_3_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_7 = T_26182_4_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_7 = T_26182_5_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_7 = T_26182_6_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_7 = T_26182_7_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_7 = T_26182_8_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_7 = T_26182_9_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_7 = T_26182_10_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_7 = T_26182_11_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_7 = T_26182_12_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_7 = T_26182_13_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_7 = T_26182_14_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_7 = T_26182_15_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_7 = T_26182_16_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_7 = T_26182_17_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_7 = T_26182_18_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_7 = T_26182_19_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_7 = T_26182_20_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_7 = T_26182_21_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_7 = T_26182_22_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_7 = T_26182_23_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_7 = T_26182_0_inst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_8 = T_26182_1_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_8 = T_26182_2_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_8 = T_26182_3_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_8 = T_26182_4_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_8 = T_26182_5_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_8 = T_26182_6_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_8 = T_26182_7_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_8 = T_26182_8_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_8 = T_26182_9_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_8 = T_26182_10_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_8 = T_26182_11_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_8 = T_26182_12_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_8 = T_26182_13_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_8 = T_26182_14_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_8 = T_26182_15_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_8 = T_26182_16_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_8 = T_26182_17_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_8 = T_26182_18_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_8 = T_26182_19_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_8 = T_26182_20_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_8 = T_26182_21_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_8 = T_26182_22_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_8 = T_26182_23_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_8 = T_26182_0_pc;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_9 = T_26182_1_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_9 = T_26182_2_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_9 = T_26182_3_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_9 = T_26182_4_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_9 = T_26182_5_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_9 = T_26182_6_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_9 = T_26182_7_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_9 = T_26182_8_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_9 = T_26182_9_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_9 = T_26182_10_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_9 = T_26182_11_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_9 = T_26182_12_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_9 = T_26182_13_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_9 = T_26182_14_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_9 = T_26182_15_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_9 = T_26182_16_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_9 = T_26182_17_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_9 = T_26182_18_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_9 = T_26182_19_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_9 = T_26182_20_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_9 = T_26182_21_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_9 = T_26182_22_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_9 = T_26182_23_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_9 = T_26182_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_10 = T_26182_1_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_10 = T_26182_2_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_10 = T_26182_3_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_10 = T_26182_4_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_10 = T_26182_5_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_10 = T_26182_6_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_10 = T_26182_7_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_10 = T_26182_8_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_10 = T_26182_9_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_10 = T_26182_10_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_10 = T_26182_11_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_10 = T_26182_12_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_10 = T_26182_13_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_10 = T_26182_14_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_10 = T_26182_15_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_10 = T_26182_16_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_10 = T_26182_17_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_10 = T_26182_18_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_10 = T_26182_19_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_10 = T_26182_20_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_10 = T_26182_21_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_10 = T_26182_22_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_10 = T_26182_23_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_10 = T_26182_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_11 = T_26182_1_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_11 = T_26182_2_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_11 = T_26182_3_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_11 = T_26182_4_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_11 = T_26182_5_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_11 = T_26182_6_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_11 = T_26182_7_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_11 = T_26182_8_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_11 = T_26182_9_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_11 = T_26182_10_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_11 = T_26182_11_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_11 = T_26182_12_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_11 = T_26182_13_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_11 = T_26182_14_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_11 = T_26182_15_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_11 = T_26182_16_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_11 = T_26182_17_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_11 = T_26182_18_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_11 = T_26182_19_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_11 = T_26182_20_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_11 = T_26182_21_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_11 = T_26182_22_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_11 = T_26182_23_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_11 = T_26182_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_12 = T_26182_1_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_12 = T_26182_2_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_12 = T_26182_3_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_12 = T_26182_4_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_12 = T_26182_5_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_12 = T_26182_6_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_12 = T_26182_7_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_12 = T_26182_8_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_12 = T_26182_9_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_12 = T_26182_10_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_12 = T_26182_11_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_12 = T_26182_12_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_12 = T_26182_13_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_12 = T_26182_14_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_12 = T_26182_15_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_12 = T_26182_16_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_12 = T_26182_17_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_12 = T_26182_18_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_12 = T_26182_19_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_12 = T_26182_20_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_12 = T_26182_21_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_12 = T_26182_22_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_12 = T_26182_23_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_12 = T_26182_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_13 = T_26182_1_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_13 = T_26182_2_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_13 = T_26182_3_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_13 = T_26182_4_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_13 = T_26182_5_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_13 = T_26182_6_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_13 = T_26182_7_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_13 = T_26182_8_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_13 = T_26182_9_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_13 = T_26182_10_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_13 = T_26182_11_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_13 = T_26182_12_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_13 = T_26182_13_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_13 = T_26182_14_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_13 = T_26182_15_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_13 = T_26182_16_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_13 = T_26182_17_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_13 = T_26182_18_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_13 = T_26182_19_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_13 = T_26182_20_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_13 = T_26182_21_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_13 = T_26182_22_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_13 = T_26182_23_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_13 = T_26182_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_14 = T_26182_1_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_14 = T_26182_2_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_14 = T_26182_3_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_14 = T_26182_4_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_14 = T_26182_5_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_14 = T_26182_6_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_14 = T_26182_7_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_14 = T_26182_8_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_14 = T_26182_9_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_14 = T_26182_10_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_14 = T_26182_11_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_14 = T_26182_12_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_14 = T_26182_13_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_14 = T_26182_14_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_14 = T_26182_15_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_14 = T_26182_16_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_14 = T_26182_17_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_14 = T_26182_18_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_14 = T_26182_19_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_14 = T_26182_20_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_14 = T_26182_21_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_14 = T_26182_22_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_14 = T_26182_23_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_14 = T_26182_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_15 = T_26182_1_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_15 = T_26182_2_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_15 = T_26182_3_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_15 = T_26182_4_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_15 = T_26182_5_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_15 = T_26182_6_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_15 = T_26182_7_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_15 = T_26182_8_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_15 = T_26182_9_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_15 = T_26182_10_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_15 = T_26182_11_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_15 = T_26182_12_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_15 = T_26182_13_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_15 = T_26182_14_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_15 = T_26182_15_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_15 = T_26182_16_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_15 = T_26182_17_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_15 = T_26182_18_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_15 = T_26182_19_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_15 = T_26182_20_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_15 = T_26182_21_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_15 = T_26182_22_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_15 = T_26182_23_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_15 = T_26182_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_16 = T_26182_1_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_16 = T_26182_2_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_16 = T_26182_3_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_16 = T_26182_4_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_16 = T_26182_5_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_16 = T_26182_6_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_16 = T_26182_7_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_16 = T_26182_8_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_16 = T_26182_9_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_16 = T_26182_10_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_16 = T_26182_11_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_16 = T_26182_12_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_16 = T_26182_13_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_16 = T_26182_14_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_16 = T_26182_15_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_16 = T_26182_16_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_16 = T_26182_17_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_16 = T_26182_18_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_16 = T_26182_19_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_16 = T_26182_20_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_16 = T_26182_21_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_16 = T_26182_22_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_16 = T_26182_23_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_16 = T_26182_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_17 = T_26182_1_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_17 = T_26182_2_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_17 = T_26182_3_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_17 = T_26182_4_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_17 = T_26182_5_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_17 = T_26182_6_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_17 = T_26182_7_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_17 = T_26182_8_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_17 = T_26182_9_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_17 = T_26182_10_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_17 = T_26182_11_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_17 = T_26182_12_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_17 = T_26182_13_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_17 = T_26182_14_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_17 = T_26182_15_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_17 = T_26182_16_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_17 = T_26182_17_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_17 = T_26182_18_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_17 = T_26182_19_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_17 = T_26182_20_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_17 = T_26182_21_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_17 = T_26182_22_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_17 = T_26182_23_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_17 = T_26182_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_18 = T_26182_1_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_18 = T_26182_2_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_18 = T_26182_3_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_18 = T_26182_4_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_18 = T_26182_5_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_18 = T_26182_6_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_18 = T_26182_7_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_18 = T_26182_8_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_18 = T_26182_9_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_18 = T_26182_10_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_18 = T_26182_11_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_18 = T_26182_12_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_18 = T_26182_13_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_18 = T_26182_14_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_18 = T_26182_15_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_18 = T_26182_16_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_18 = T_26182_17_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_18 = T_26182_18_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_18 = T_26182_19_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_18 = T_26182_20_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_18 = T_26182_21_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_18 = T_26182_22_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_18 = T_26182_23_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_18 = T_26182_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_19 = T_26182_1_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_19 = T_26182_2_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_19 = T_26182_3_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_19 = T_26182_4_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_19 = T_26182_5_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_19 = T_26182_6_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_19 = T_26182_7_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_19 = T_26182_8_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_19 = T_26182_9_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_19 = T_26182_10_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_19 = T_26182_11_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_19 = T_26182_12_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_19 = T_26182_13_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_19 = T_26182_14_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_19 = T_26182_15_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_19 = T_26182_16_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_19 = T_26182_17_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_19 = T_26182_18_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_19 = T_26182_19_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_19 = T_26182_20_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_19 = T_26182_21_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_19 = T_26182_22_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_19 = T_26182_23_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_19 = T_26182_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_20 = T_26182_1_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_20 = T_26182_2_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_20 = T_26182_3_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_20 = T_26182_4_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_20 = T_26182_5_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_20 = T_26182_6_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_20 = T_26182_7_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_20 = T_26182_8_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_20 = T_26182_9_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_20 = T_26182_10_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_20 = T_26182_11_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_20 = T_26182_12_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_20 = T_26182_13_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_20 = T_26182_14_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_20 = T_26182_15_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_20 = T_26182_16_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_20 = T_26182_17_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_20 = T_26182_18_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_20 = T_26182_19_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_20 = T_26182_20_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_20 = T_26182_21_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_20 = T_26182_22_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_20 = T_26182_23_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_20 = T_26182_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_21 = T_26182_1_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_21 = T_26182_2_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_21 = T_26182_3_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_21 = T_26182_4_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_21 = T_26182_5_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_21 = T_26182_6_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_21 = T_26182_7_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_21 = T_26182_8_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_21 = T_26182_9_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_21 = T_26182_10_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_21 = T_26182_11_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_21 = T_26182_12_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_21 = T_26182_13_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_21 = T_26182_14_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_21 = T_26182_15_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_21 = T_26182_16_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_21 = T_26182_17_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_21 = T_26182_18_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_21 = T_26182_19_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_21 = T_26182_20_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_21 = T_26182_21_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_21 = T_26182_22_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_21 = T_26182_23_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_21 = T_26182_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_22 = T_26182_1_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_22 = T_26182_2_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_22 = T_26182_3_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_22 = T_26182_4_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_22 = T_26182_5_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_22 = T_26182_6_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_22 = T_26182_7_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_22 = T_26182_8_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_22 = T_26182_9_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_22 = T_26182_10_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_22 = T_26182_11_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_22 = T_26182_12_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_22 = T_26182_13_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_22 = T_26182_14_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_22 = T_26182_15_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_22 = T_26182_16_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_22 = T_26182_17_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_22 = T_26182_18_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_22 = T_26182_19_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_22 = T_26182_20_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_22 = T_26182_21_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_22 = T_26182_22_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_22 = T_26182_23_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_22 = T_26182_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_23 = T_26182_1_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_23 = T_26182_2_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_23 = T_26182_3_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_23 = T_26182_4_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_23 = T_26182_5_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_23 = T_26182_6_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_23 = T_26182_7_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_23 = T_26182_8_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_23 = T_26182_9_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_23 = T_26182_10_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_23 = T_26182_11_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_23 = T_26182_12_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_23 = T_26182_13_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_23 = T_26182_14_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_23 = T_26182_15_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_23 = T_26182_16_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_23 = T_26182_17_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_23 = T_26182_18_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_23 = T_26182_19_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_23 = T_26182_20_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_23 = T_26182_21_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_23 = T_26182_22_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_23 = T_26182_23_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_23 = T_26182_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_24 = T_26182_1_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_24 = T_26182_2_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_24 = T_26182_3_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_24 = T_26182_4_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_24 = T_26182_5_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_24 = T_26182_6_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_24 = T_26182_7_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_24 = T_26182_8_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_24 = T_26182_9_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_24 = T_26182_10_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_24 = T_26182_11_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_24 = T_26182_12_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_24 = T_26182_13_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_24 = T_26182_14_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_24 = T_26182_15_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_24 = T_26182_16_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_24 = T_26182_17_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_24 = T_26182_18_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_24 = T_26182_19_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_24 = T_26182_20_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_24 = T_26182_21_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_24 = T_26182_22_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_24 = T_26182_23_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_24 = T_26182_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_25 = T_26182_1_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_25 = T_26182_2_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_25 = T_26182_3_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_25 = T_26182_4_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_25 = T_26182_5_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_25 = T_26182_6_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_25 = T_26182_7_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_25 = T_26182_8_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_25 = T_26182_9_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_25 = T_26182_10_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_25 = T_26182_11_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_25 = T_26182_12_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_25 = T_26182_13_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_25 = T_26182_14_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_25 = T_26182_15_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_25 = T_26182_16_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_25 = T_26182_17_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_25 = T_26182_18_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_25 = T_26182_19_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_25 = T_26182_20_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_25 = T_26182_21_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_25 = T_26182_22_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_25 = T_26182_23_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_25 = T_26182_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_26 = T_26182_1_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_26 = T_26182_2_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_26 = T_26182_3_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_26 = T_26182_4_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_26 = T_26182_5_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_26 = T_26182_6_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_26 = T_26182_7_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_26 = T_26182_8_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_26 = T_26182_9_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_26 = T_26182_10_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_26 = T_26182_11_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_26 = T_26182_12_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_26 = T_26182_13_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_26 = T_26182_14_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_26 = T_26182_15_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_26 = T_26182_16_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_26 = T_26182_17_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_26 = T_26182_18_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_26 = T_26182_19_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_26 = T_26182_20_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_26 = T_26182_21_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_26 = T_26182_22_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_26 = T_26182_23_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_26 = T_26182_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_27 = T_26182_1_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_27 = T_26182_2_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_27 = T_26182_3_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_27 = T_26182_4_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_27 = T_26182_5_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_27 = T_26182_6_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_27 = T_26182_7_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_27 = T_26182_8_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_27 = T_26182_9_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_27 = T_26182_10_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_27 = T_26182_11_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_27 = T_26182_12_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_27 = T_26182_13_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_27 = T_26182_14_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_27 = T_26182_15_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_27 = T_26182_16_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_27 = T_26182_17_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_27 = T_26182_18_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_27 = T_26182_19_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_27 = T_26182_20_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_27 = T_26182_21_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_27 = T_26182_22_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_27 = T_26182_23_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_27 = T_26182_0_is_call;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_28 = T_26182_1_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_28 = T_26182_2_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_28 = T_26182_3_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_28 = T_26182_4_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_28 = T_26182_5_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_28 = T_26182_6_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_28 = T_26182_7_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_28 = T_26182_8_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_28 = T_26182_9_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_28 = T_26182_10_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_28 = T_26182_11_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_28 = T_26182_12_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_28 = T_26182_13_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_28 = T_26182_14_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_28 = T_26182_15_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_28 = T_26182_16_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_28 = T_26182_17_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_28 = T_26182_18_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_28 = T_26182_19_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_28 = T_26182_20_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_28 = T_26182_21_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_28 = T_26182_22_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_28 = T_26182_23_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_28 = T_26182_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_29 = T_26182_1_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_29 = T_26182_2_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_29 = T_26182_3_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_29 = T_26182_4_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_29 = T_26182_5_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_29 = T_26182_6_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_29 = T_26182_7_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_29 = T_26182_8_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_29 = T_26182_9_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_29 = T_26182_10_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_29 = T_26182_11_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_29 = T_26182_12_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_29 = T_26182_13_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_29 = T_26182_14_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_29 = T_26182_15_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_29 = T_26182_16_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_29 = T_26182_17_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_29 = T_26182_18_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_29 = T_26182_19_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_29 = T_26182_20_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_29 = T_26182_21_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_29 = T_26182_22_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_29 = T_26182_23_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_29 = T_26182_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_30 = T_26182_1_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_30 = T_26182_2_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_30 = T_26182_3_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_30 = T_26182_4_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_30 = T_26182_5_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_30 = T_26182_6_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_30 = T_26182_7_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_30 = T_26182_8_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_30 = T_26182_9_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_30 = T_26182_10_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_30 = T_26182_11_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_30 = T_26182_12_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_30 = T_26182_13_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_30 = T_26182_14_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_30 = T_26182_15_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_30 = T_26182_16_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_30 = T_26182_17_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_30 = T_26182_18_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_30 = T_26182_19_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_30 = T_26182_20_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_30 = T_26182_21_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_30 = T_26182_22_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_30 = T_26182_23_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_30 = T_26182_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_31 = T_26182_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_31 = T_26182_2_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_31 = T_26182_3_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_31 = T_26182_4_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_31 = T_26182_5_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_31 = T_26182_6_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_31 = T_26182_7_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_31 = T_26182_8_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_31 = T_26182_9_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_31 = T_26182_10_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_31 = T_26182_11_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_31 = T_26182_12_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_31 = T_26182_13_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_31 = T_26182_14_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_31 = T_26182_15_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_31 = T_26182_16_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_31 = T_26182_17_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_31 = T_26182_18_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_31 = T_26182_19_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_31 = T_26182_20_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_31 = T_26182_21_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_31 = T_26182_22_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_31 = T_26182_23_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_31 = T_26182_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_32 = T_26182_1_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_32 = T_26182_2_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_32 = T_26182_3_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_32 = T_26182_4_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_32 = T_26182_5_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_32 = T_26182_6_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_32 = T_26182_7_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_32 = T_26182_8_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_32 = T_26182_9_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_32 = T_26182_10_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_32 = T_26182_11_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_32 = T_26182_12_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_32 = T_26182_13_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_32 = T_26182_14_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_32 = T_26182_15_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_32 = T_26182_16_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_32 = T_26182_17_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_32 = T_26182_18_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_32 = T_26182_19_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_32 = T_26182_20_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_32 = T_26182_21_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_32 = T_26182_22_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_32 = T_26182_23_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_32 = T_26182_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_33 = T_26182_1_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_33 = T_26182_2_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_33 = T_26182_3_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_33 = T_26182_4_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_33 = T_26182_5_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_33 = T_26182_6_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_33 = T_26182_7_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_33 = T_26182_8_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_33 = T_26182_9_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_33 = T_26182_10_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_33 = T_26182_11_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_33 = T_26182_12_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_33 = T_26182_13_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_33 = T_26182_14_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_33 = T_26182_15_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_33 = T_26182_16_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_33 = T_26182_17_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_33 = T_26182_18_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_33 = T_26182_19_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_33 = T_26182_20_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_33 = T_26182_21_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_33 = T_26182_22_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_33 = T_26182_23_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_33 = T_26182_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_34 = T_26182_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_34 = T_26182_2_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_34 = T_26182_3_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_34 = T_26182_4_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_34 = T_26182_5_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_34 = T_26182_6_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_34 = T_26182_7_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_34 = T_26182_8_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_34 = T_26182_9_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_34 = T_26182_10_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_34 = T_26182_11_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_34 = T_26182_12_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_34 = T_26182_13_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_34 = T_26182_14_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_34 = T_26182_15_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_34 = T_26182_16_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_34 = T_26182_17_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_34 = T_26182_18_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_34 = T_26182_19_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_34 = T_26182_20_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_34 = T_26182_21_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_34 = T_26182_22_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_34 = T_26182_23_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_34 = T_26182_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_35 = T_26182_1_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_35 = T_26182_2_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_35 = T_26182_3_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_35 = T_26182_4_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_35 = T_26182_5_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_35 = T_26182_6_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_35 = T_26182_7_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_35 = T_26182_8_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_35 = T_26182_9_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_35 = T_26182_10_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_35 = T_26182_11_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_35 = T_26182_12_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_35 = T_26182_13_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_35 = T_26182_14_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_35 = T_26182_15_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_35 = T_26182_16_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_35 = T_26182_17_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_35 = T_26182_18_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_35 = T_26182_19_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_35 = T_26182_20_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_35 = T_26182_21_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_35 = T_26182_22_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_35 = T_26182_23_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_35 = T_26182_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_36 = T_26182_1_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_36 = T_26182_2_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_36 = T_26182_3_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_36 = T_26182_4_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_36 = T_26182_5_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_36 = T_26182_6_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_36 = T_26182_7_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_36 = T_26182_8_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_36 = T_26182_9_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_36 = T_26182_10_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_36 = T_26182_11_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_36 = T_26182_12_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_36 = T_26182_13_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_36 = T_26182_14_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_36 = T_26182_15_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_36 = T_26182_16_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_36 = T_26182_17_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_36 = T_26182_18_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_36 = T_26182_19_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_36 = T_26182_20_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_36 = T_26182_21_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_36 = T_26182_22_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_36 = T_26182_23_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_36 = T_26182_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_37 = T_26182_1_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_37 = T_26182_2_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_37 = T_26182_3_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_37 = T_26182_4_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_37 = T_26182_5_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_37 = T_26182_6_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_37 = T_26182_7_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_37 = T_26182_8_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_37 = T_26182_9_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_37 = T_26182_10_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_37 = T_26182_11_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_37 = T_26182_12_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_37 = T_26182_13_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_37 = T_26182_14_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_37 = T_26182_15_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_37 = T_26182_16_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_37 = T_26182_17_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_37 = T_26182_18_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_37 = T_26182_19_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_37 = T_26182_20_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_37 = T_26182_21_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_37 = T_26182_22_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_37 = T_26182_23_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_37 = T_26182_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_38 = T_26182_1_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_38 = T_26182_2_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_38 = T_26182_3_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_38 = T_26182_4_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_38 = T_26182_5_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_38 = T_26182_6_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_38 = T_26182_7_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_38 = T_26182_8_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_38 = T_26182_9_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_38 = T_26182_10_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_38 = T_26182_11_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_38 = T_26182_12_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_38 = T_26182_13_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_38 = T_26182_14_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_38 = T_26182_15_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_38 = T_26182_16_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_38 = T_26182_17_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_38 = T_26182_18_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_38 = T_26182_19_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_38 = T_26182_20_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_38 = T_26182_21_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_38 = T_26182_22_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_38 = T_26182_23_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_38 = T_26182_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_39 = T_26182_1_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_39 = T_26182_2_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_39 = T_26182_3_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_39 = T_26182_4_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_39 = T_26182_5_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_39 = T_26182_6_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_39 = T_26182_7_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_39 = T_26182_8_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_39 = T_26182_9_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_39 = T_26182_10_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_39 = T_26182_11_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_39 = T_26182_12_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_39 = T_26182_13_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_39 = T_26182_14_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_39 = T_26182_15_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_39 = T_26182_16_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_39 = T_26182_17_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_39 = T_26182_18_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_39 = T_26182_19_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_39 = T_26182_20_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_39 = T_26182_21_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_39 = T_26182_22_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_39 = T_26182_23_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_39 = T_26182_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_40 = T_26182_1_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_40 = T_26182_2_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_40 = T_26182_3_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_40 = T_26182_4_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_40 = T_26182_5_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_40 = T_26182_6_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_40 = T_26182_7_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_40 = T_26182_8_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_40 = T_26182_9_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_40 = T_26182_10_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_40 = T_26182_11_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_40 = T_26182_12_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_40 = T_26182_13_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_40 = T_26182_14_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_40 = T_26182_15_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_40 = T_26182_16_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_40 = T_26182_17_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_40 = T_26182_18_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_40 = T_26182_19_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_40 = T_26182_20_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_40 = T_26182_21_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_40 = T_26182_22_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_40 = T_26182_23_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_40 = T_26182_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_41 = T_26182_1_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_41 = T_26182_2_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_41 = T_26182_3_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_41 = T_26182_4_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_41 = T_26182_5_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_41 = T_26182_6_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_41 = T_26182_7_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_41 = T_26182_8_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_41 = T_26182_9_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_41 = T_26182_10_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_41 = T_26182_11_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_41 = T_26182_12_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_41 = T_26182_13_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_41 = T_26182_14_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_41 = T_26182_15_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_41 = T_26182_16_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_41 = T_26182_17_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_41 = T_26182_18_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_41 = T_26182_19_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_41 = T_26182_20_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_41 = T_26182_21_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_41 = T_26182_22_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_41 = T_26182_23_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_41 = T_26182_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_42 = T_26182_1_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_42 = T_26182_2_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_42 = T_26182_3_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_42 = T_26182_4_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_42 = T_26182_5_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_42 = T_26182_6_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_42 = T_26182_7_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_42 = T_26182_8_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_42 = T_26182_9_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_42 = T_26182_10_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_42 = T_26182_11_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_42 = T_26182_12_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_42 = T_26182_13_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_42 = T_26182_14_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_42 = T_26182_15_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_42 = T_26182_16_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_42 = T_26182_17_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_42 = T_26182_18_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_42 = T_26182_19_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_42 = T_26182_20_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_42 = T_26182_21_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_42 = T_26182_22_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_42 = T_26182_23_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_42 = T_26182_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_43 = T_26182_1_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_43 = T_26182_2_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_43 = T_26182_3_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_43 = T_26182_4_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_43 = T_26182_5_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_43 = T_26182_6_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_43 = T_26182_7_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_43 = T_26182_8_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_43 = T_26182_9_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_43 = T_26182_10_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_43 = T_26182_11_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_43 = T_26182_12_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_43 = T_26182_13_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_43 = T_26182_14_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_43 = T_26182_15_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_43 = T_26182_16_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_43 = T_26182_17_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_43 = T_26182_18_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_43 = T_26182_19_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_43 = T_26182_20_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_43 = T_26182_21_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_43 = T_26182_22_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_43 = T_26182_23_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_43 = T_26182_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_44 = T_26182_1_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_44 = T_26182_2_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_44 = T_26182_3_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_44 = T_26182_4_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_44 = T_26182_5_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_44 = T_26182_6_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_44 = T_26182_7_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_44 = T_26182_8_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_44 = T_26182_9_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_44 = T_26182_10_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_44 = T_26182_11_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_44 = T_26182_12_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_44 = T_26182_13_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_44 = T_26182_14_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_44 = T_26182_15_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_44 = T_26182_16_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_44 = T_26182_17_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_44 = T_26182_18_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_44 = T_26182_19_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_44 = T_26182_20_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_44 = T_26182_21_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_44 = T_26182_22_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_44 = T_26182_23_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_44 = T_26182_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_45 = T_26182_1_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_45 = T_26182_2_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_45 = T_26182_3_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_45 = T_26182_4_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_45 = T_26182_5_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_45 = T_26182_6_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_45 = T_26182_7_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_45 = T_26182_8_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_45 = T_26182_9_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_45 = T_26182_10_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_45 = T_26182_11_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_45 = T_26182_12_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_45 = T_26182_13_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_45 = T_26182_14_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_45 = T_26182_15_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_45 = T_26182_16_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_45 = T_26182_17_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_45 = T_26182_18_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_45 = T_26182_19_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_45 = T_26182_20_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_45 = T_26182_21_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_45 = T_26182_22_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_45 = T_26182_23_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_45 = T_26182_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_46 = T_26182_1_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_46 = T_26182_2_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_46 = T_26182_3_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_46 = T_26182_4_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_46 = T_26182_5_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_46 = T_26182_6_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_46 = T_26182_7_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_46 = T_26182_8_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_46 = T_26182_9_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_46 = T_26182_10_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_46 = T_26182_11_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_46 = T_26182_12_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_46 = T_26182_13_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_46 = T_26182_14_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_46 = T_26182_15_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_46 = T_26182_16_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_46 = T_26182_17_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_46 = T_26182_18_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_46 = T_26182_19_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_46 = T_26182_20_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_46 = T_26182_21_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_46 = T_26182_22_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_46 = T_26182_23_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_46 = T_26182_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_47 = T_26182_1_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_47 = T_26182_2_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_47 = T_26182_3_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_47 = T_26182_4_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_47 = T_26182_5_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_47 = T_26182_6_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_47 = T_26182_7_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_47 = T_26182_8_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_47 = T_26182_9_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_47 = T_26182_10_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_47 = T_26182_11_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_47 = T_26182_12_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_47 = T_26182_13_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_47 = T_26182_14_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_47 = T_26182_15_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_47 = T_26182_16_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_47 = T_26182_17_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_47 = T_26182_18_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_47 = T_26182_19_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_47 = T_26182_20_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_47 = T_26182_21_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_47 = T_26182_22_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_47 = T_26182_23_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_47 = T_26182_0_pdst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_48 = T_26182_1_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_48 = T_26182_2_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_48 = T_26182_3_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_48 = T_26182_4_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_48 = T_26182_5_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_48 = T_26182_6_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_48 = T_26182_7_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_48 = T_26182_8_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_48 = T_26182_9_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_48 = T_26182_10_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_48 = T_26182_11_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_48 = T_26182_12_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_48 = T_26182_13_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_48 = T_26182_14_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_48 = T_26182_15_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_48 = T_26182_16_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_48 = T_26182_17_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_48 = T_26182_18_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_48 = T_26182_19_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_48 = T_26182_20_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_48 = T_26182_21_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_48 = T_26182_22_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_48 = T_26182_23_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_48 = T_26182_0_pop1;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_49 = T_26182_1_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_49 = T_26182_2_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_49 = T_26182_3_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_49 = T_26182_4_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_49 = T_26182_5_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_49 = T_26182_6_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_49 = T_26182_7_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_49 = T_26182_8_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_49 = T_26182_9_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_49 = T_26182_10_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_49 = T_26182_11_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_49 = T_26182_12_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_49 = T_26182_13_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_49 = T_26182_14_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_49 = T_26182_15_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_49 = T_26182_16_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_49 = T_26182_17_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_49 = T_26182_18_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_49 = T_26182_19_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_49 = T_26182_20_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_49 = T_26182_21_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_49 = T_26182_22_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_49 = T_26182_23_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_49 = T_26182_0_pop2;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_50 = T_26182_1_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_50 = T_26182_2_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_50 = T_26182_3_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_50 = T_26182_4_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_50 = T_26182_5_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_50 = T_26182_6_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_50 = T_26182_7_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_50 = T_26182_8_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_50 = T_26182_9_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_50 = T_26182_10_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_50 = T_26182_11_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_50 = T_26182_12_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_50 = T_26182_13_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_50 = T_26182_14_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_50 = T_26182_15_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_50 = T_26182_16_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_50 = T_26182_17_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_50 = T_26182_18_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_50 = T_26182_19_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_50 = T_26182_20_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_50 = T_26182_21_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_50 = T_26182_22_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_50 = T_26182_23_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_50 = T_26182_0_pop3;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_51 = T_26182_1_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_51 = T_26182_2_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_51 = T_26182_3_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_51 = T_26182_4_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_51 = T_26182_5_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_51 = T_26182_6_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_51 = T_26182_7_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_51 = T_26182_8_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_51 = T_26182_9_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_51 = T_26182_10_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_51 = T_26182_11_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_51 = T_26182_12_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_51 = T_26182_13_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_51 = T_26182_14_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_51 = T_26182_15_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_51 = T_26182_16_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_51 = T_26182_17_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_51 = T_26182_18_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_51 = T_26182_19_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_51 = T_26182_20_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_51 = T_26182_21_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_51 = T_26182_22_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_51 = T_26182_23_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_51 = T_26182_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_52 = T_26182_1_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_52 = T_26182_2_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_52 = T_26182_3_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_52 = T_26182_4_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_52 = T_26182_5_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_52 = T_26182_6_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_52 = T_26182_7_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_52 = T_26182_8_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_52 = T_26182_9_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_52 = T_26182_10_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_52 = T_26182_11_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_52 = T_26182_12_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_52 = T_26182_13_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_52 = T_26182_14_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_52 = T_26182_15_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_52 = T_26182_16_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_52 = T_26182_17_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_52 = T_26182_18_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_52 = T_26182_19_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_52 = T_26182_20_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_52 = T_26182_21_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_52 = T_26182_22_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_52 = T_26182_23_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_52 = T_26182_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_53 = T_26182_1_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_53 = T_26182_2_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_53 = T_26182_3_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_53 = T_26182_4_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_53 = T_26182_5_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_53 = T_26182_6_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_53 = T_26182_7_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_53 = T_26182_8_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_53 = T_26182_9_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_53 = T_26182_10_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_53 = T_26182_11_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_53 = T_26182_12_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_53 = T_26182_13_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_53 = T_26182_14_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_53 = T_26182_15_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_53 = T_26182_16_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_53 = T_26182_17_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_53 = T_26182_18_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_53 = T_26182_19_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_53 = T_26182_20_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_53 = T_26182_21_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_53 = T_26182_22_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_53 = T_26182_23_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_53 = T_26182_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_54 = T_26182_1_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_54 = T_26182_2_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_54 = T_26182_3_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_54 = T_26182_4_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_54 = T_26182_5_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_54 = T_26182_6_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_54 = T_26182_7_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_54 = T_26182_8_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_54 = T_26182_9_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_54 = T_26182_10_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_54 = T_26182_11_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_54 = T_26182_12_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_54 = T_26182_13_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_54 = T_26182_14_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_54 = T_26182_15_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_54 = T_26182_16_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_54 = T_26182_17_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_54 = T_26182_18_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_54 = T_26182_19_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_54 = T_26182_20_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_54 = T_26182_21_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_54 = T_26182_22_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_54 = T_26182_23_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_54 = T_26182_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_55 = T_26182_1_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_55 = T_26182_2_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_55 = T_26182_3_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_55 = T_26182_4_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_55 = T_26182_5_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_55 = T_26182_6_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_55 = T_26182_7_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_55 = T_26182_8_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_55 = T_26182_9_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_55 = T_26182_10_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_55 = T_26182_11_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_55 = T_26182_12_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_55 = T_26182_13_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_55 = T_26182_14_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_55 = T_26182_15_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_55 = T_26182_16_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_55 = T_26182_17_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_55 = T_26182_18_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_55 = T_26182_19_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_55 = T_26182_20_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_55 = T_26182_21_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_55 = T_26182_22_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_55 = T_26182_23_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_55 = T_26182_0_exception;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_56 = T_26182_1_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_56 = T_26182_2_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_56 = T_26182_3_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_56 = T_26182_4_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_56 = T_26182_5_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_56 = T_26182_6_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_56 = T_26182_7_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_56 = T_26182_8_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_56 = T_26182_9_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_56 = T_26182_10_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_56 = T_26182_11_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_56 = T_26182_12_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_56 = T_26182_13_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_56 = T_26182_14_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_56 = T_26182_15_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_56 = T_26182_16_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_56 = T_26182_17_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_56 = T_26182_18_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_56 = T_26182_19_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_56 = T_26182_20_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_56 = T_26182_21_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_56 = T_26182_22_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_56 = T_26182_23_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_56 = T_26182_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_57 = T_26182_1_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_57 = T_26182_2_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_57 = T_26182_3_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_57 = T_26182_4_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_57 = T_26182_5_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_57 = T_26182_6_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_57 = T_26182_7_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_57 = T_26182_8_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_57 = T_26182_9_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_57 = T_26182_10_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_57 = T_26182_11_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_57 = T_26182_12_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_57 = T_26182_13_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_57 = T_26182_14_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_57 = T_26182_15_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_57 = T_26182_16_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_57 = T_26182_17_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_57 = T_26182_18_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_57 = T_26182_19_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_57 = T_26182_20_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_57 = T_26182_21_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_57 = T_26182_22_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_57 = T_26182_23_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_57 = T_26182_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_58 = T_26182_1_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_58 = T_26182_2_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_58 = T_26182_3_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_58 = T_26182_4_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_58 = T_26182_5_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_58 = T_26182_6_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_58 = T_26182_7_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_58 = T_26182_8_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_58 = T_26182_9_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_58 = T_26182_10_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_58 = T_26182_11_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_58 = T_26182_12_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_58 = T_26182_13_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_58 = T_26182_14_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_58 = T_26182_15_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_58 = T_26182_16_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_58 = T_26182_17_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_58 = T_26182_18_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_58 = T_26182_19_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_58 = T_26182_20_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_58 = T_26182_21_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_58 = T_26182_22_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_58 = T_26182_23_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_58 = T_26182_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_59 = T_26182_1_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_59 = T_26182_2_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_59 = T_26182_3_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_59 = T_26182_4_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_59 = T_26182_5_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_59 = T_26182_6_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_59 = T_26182_7_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_59 = T_26182_8_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_59 = T_26182_9_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_59 = T_26182_10_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_59 = T_26182_11_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_59 = T_26182_12_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_59 = T_26182_13_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_59 = T_26182_14_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_59 = T_26182_15_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_59 = T_26182_16_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_59 = T_26182_17_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_59 = T_26182_18_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_59 = T_26182_19_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_59 = T_26182_20_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_59 = T_26182_21_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_59 = T_26182_22_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_59 = T_26182_23_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_59 = T_26182_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_60 = T_26182_1_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_60 = T_26182_2_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_60 = T_26182_3_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_60 = T_26182_4_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_60 = T_26182_5_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_60 = T_26182_6_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_60 = T_26182_7_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_60 = T_26182_8_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_60 = T_26182_9_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_60 = T_26182_10_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_60 = T_26182_11_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_60 = T_26182_12_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_60 = T_26182_13_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_60 = T_26182_14_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_60 = T_26182_15_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_60 = T_26182_16_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_60 = T_26182_17_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_60 = T_26182_18_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_60 = T_26182_19_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_60 = T_26182_20_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_60 = T_26182_21_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_60 = T_26182_22_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_60 = T_26182_23_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_60 = T_26182_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_61 = T_26182_1_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_61 = T_26182_2_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_61 = T_26182_3_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_61 = T_26182_4_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_61 = T_26182_5_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_61 = T_26182_6_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_61 = T_26182_7_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_61 = T_26182_8_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_61 = T_26182_9_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_61 = T_26182_10_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_61 = T_26182_11_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_61 = T_26182_12_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_61 = T_26182_13_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_61 = T_26182_14_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_61 = T_26182_15_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_61 = T_26182_16_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_61 = T_26182_17_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_61 = T_26182_18_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_61 = T_26182_19_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_61 = T_26182_20_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_61 = T_26182_21_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_61 = T_26182_22_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_61 = T_26182_23_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_61 = T_26182_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_62 = T_26182_1_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_62 = T_26182_2_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_62 = T_26182_3_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_62 = T_26182_4_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_62 = T_26182_5_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_62 = T_26182_6_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_62 = T_26182_7_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_62 = T_26182_8_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_62 = T_26182_9_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_62 = T_26182_10_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_62 = T_26182_11_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_62 = T_26182_12_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_62 = T_26182_13_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_62 = T_26182_14_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_62 = T_26182_15_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_62 = T_26182_16_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_62 = T_26182_17_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_62 = T_26182_18_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_62 = T_26182_19_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_62 = T_26182_20_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_62 = T_26182_21_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_62 = T_26182_22_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_62 = T_26182_23_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_62 = T_26182_0_is_store;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_63 = T_26182_1_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_63 = T_26182_2_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_63 = T_26182_3_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_63 = T_26182_4_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_63 = T_26182_5_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_63 = T_26182_6_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_63 = T_26182_7_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_63 = T_26182_8_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_63 = T_26182_9_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_63 = T_26182_10_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_63 = T_26182_11_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_63 = T_26182_12_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_63 = T_26182_13_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_63 = T_26182_14_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_63 = T_26182_15_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_63 = T_26182_16_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_63 = T_26182_17_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_63 = T_26182_18_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_63 = T_26182_19_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_63 = T_26182_20_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_63 = T_26182_21_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_63 = T_26182_22_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_63 = T_26182_23_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_63 = T_26182_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_64 = T_26182_1_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_64 = T_26182_2_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_64 = T_26182_3_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_64 = T_26182_4_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_64 = T_26182_5_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_64 = T_26182_6_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_64 = T_26182_7_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_64 = T_26182_8_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_64 = T_26182_9_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_64 = T_26182_10_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_64 = T_26182_11_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_64 = T_26182_12_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_64 = T_26182_13_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_64 = T_26182_14_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_64 = T_26182_15_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_64 = T_26182_16_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_64 = T_26182_17_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_64 = T_26182_18_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_64 = T_26182_19_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_64 = T_26182_20_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_64 = T_26182_21_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_64 = T_26182_22_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_64 = T_26182_23_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_64 = T_26182_0_is_load;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_65 = T_26182_1_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_65 = T_26182_2_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_65 = T_26182_3_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_65 = T_26182_4_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_65 = T_26182_5_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_65 = T_26182_6_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_65 = T_26182_7_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_65 = T_26182_8_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_65 = T_26182_9_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_65 = T_26182_10_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_65 = T_26182_11_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_65 = T_26182_12_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_65 = T_26182_13_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_65 = T_26182_14_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_65 = T_26182_15_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_65 = T_26182_16_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_65 = T_26182_17_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_65 = T_26182_18_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_65 = T_26182_19_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_65 = T_26182_20_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_65 = T_26182_21_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_65 = T_26182_22_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_65 = T_26182_23_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_65 = T_26182_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_66 = T_26182_1_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_66 = T_26182_2_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_66 = T_26182_3_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_66 = T_26182_4_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_66 = T_26182_5_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_66 = T_26182_6_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_66 = T_26182_7_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_66 = T_26182_8_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_66 = T_26182_9_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_66 = T_26182_10_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_66 = T_26182_11_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_66 = T_26182_12_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_66 = T_26182_13_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_66 = T_26182_14_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_66 = T_26182_15_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_66 = T_26182_16_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_66 = T_26182_17_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_66 = T_26182_18_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_66 = T_26182_19_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_66 = T_26182_20_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_66 = T_26182_21_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_66 = T_26182_22_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_66 = T_26182_23_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_66 = T_26182_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_67 = T_26182_1_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_67 = T_26182_2_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_67 = T_26182_3_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_67 = T_26182_4_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_67 = T_26182_5_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_67 = T_26182_6_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_67 = T_26182_7_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_67 = T_26182_8_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_67 = T_26182_9_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_67 = T_26182_10_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_67 = T_26182_11_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_67 = T_26182_12_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_67 = T_26182_13_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_67 = T_26182_14_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_67 = T_26182_15_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_67 = T_26182_16_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_67 = T_26182_17_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_67 = T_26182_18_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_67 = T_26182_19_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_67 = T_26182_20_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_67 = T_26182_21_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_67 = T_26182_22_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_67 = T_26182_23_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_67 = T_26182_0_ldst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_68 = T_26182_1_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_68 = T_26182_2_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_68 = T_26182_3_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_68 = T_26182_4_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_68 = T_26182_5_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_68 = T_26182_6_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_68 = T_26182_7_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_68 = T_26182_8_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_68 = T_26182_9_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_68 = T_26182_10_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_68 = T_26182_11_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_68 = T_26182_12_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_68 = T_26182_13_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_68 = T_26182_14_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_68 = T_26182_15_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_68 = T_26182_16_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_68 = T_26182_17_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_68 = T_26182_18_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_68 = T_26182_19_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_68 = T_26182_20_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_68 = T_26182_21_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_68 = T_26182_22_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_68 = T_26182_23_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_68 = T_26182_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_69 = T_26182_1_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_69 = T_26182_2_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_69 = T_26182_3_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_69 = T_26182_4_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_69 = T_26182_5_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_69 = T_26182_6_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_69 = T_26182_7_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_69 = T_26182_8_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_69 = T_26182_9_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_69 = T_26182_10_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_69 = T_26182_11_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_69 = T_26182_12_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_69 = T_26182_13_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_69 = T_26182_14_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_69 = T_26182_15_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_69 = T_26182_16_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_69 = T_26182_17_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_69 = T_26182_18_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_69 = T_26182_19_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_69 = T_26182_20_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_69 = T_26182_21_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_69 = T_26182_22_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_69 = T_26182_23_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_69 = T_26182_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_70 = T_26182_1_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_70 = T_26182_2_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_70 = T_26182_3_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_70 = T_26182_4_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_70 = T_26182_5_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_70 = T_26182_6_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_70 = T_26182_7_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_70 = T_26182_8_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_70 = T_26182_9_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_70 = T_26182_10_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_70 = T_26182_11_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_70 = T_26182_12_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_70 = T_26182_13_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_70 = T_26182_14_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_70 = T_26182_15_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_70 = T_26182_16_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_70 = T_26182_17_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_70 = T_26182_18_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_70 = T_26182_19_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_70 = T_26182_20_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_70 = T_26182_21_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_70 = T_26182_22_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_70 = T_26182_23_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_70 = T_26182_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_71 = T_26182_1_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_71 = T_26182_2_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_71 = T_26182_3_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_71 = T_26182_4_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_71 = T_26182_5_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_71 = T_26182_6_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_71 = T_26182_7_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_71 = T_26182_8_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_71 = T_26182_9_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_71 = T_26182_10_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_71 = T_26182_11_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_71 = T_26182_12_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_71 = T_26182_13_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_71 = T_26182_14_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_71 = T_26182_15_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_71 = T_26182_16_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_71 = T_26182_17_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_71 = T_26182_18_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_71 = T_26182_19_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_71 = T_26182_20_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_71 = T_26182_21_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_71 = T_26182_22_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_71 = T_26182_23_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_71 = T_26182_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_72 = T_26182_1_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_72 = T_26182_2_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_72 = T_26182_3_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_72 = T_26182_4_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_72 = T_26182_5_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_72 = T_26182_6_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_72 = T_26182_7_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_72 = T_26182_8_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_72 = T_26182_9_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_72 = T_26182_10_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_72 = T_26182_11_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_72 = T_26182_12_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_72 = T_26182_13_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_72 = T_26182_14_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_72 = T_26182_15_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_72 = T_26182_16_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_72 = T_26182_17_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_72 = T_26182_18_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_72 = T_26182_19_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_72 = T_26182_20_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_72 = T_26182_21_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_72 = T_26182_22_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_72 = T_26182_23_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_72 = T_26182_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_73 = T_26182_1_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_73 = T_26182_2_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_73 = T_26182_3_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_73 = T_26182_4_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_73 = T_26182_5_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_73 = T_26182_6_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_73 = T_26182_7_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_73 = T_26182_8_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_73 = T_26182_9_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_73 = T_26182_10_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_73 = T_26182_11_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_73 = T_26182_12_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_73 = T_26182_13_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_73 = T_26182_14_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_73 = T_26182_15_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_73 = T_26182_16_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_73 = T_26182_17_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_73 = T_26182_18_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_73 = T_26182_19_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_73 = T_26182_20_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_73 = T_26182_21_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_73 = T_26182_22_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_73 = T_26182_23_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_73 = T_26182_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_74 = T_26182_1_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_74 = T_26182_2_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_74 = T_26182_3_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_74 = T_26182_4_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_74 = T_26182_5_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_74 = T_26182_6_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_74 = T_26182_7_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_74 = T_26182_8_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_74 = T_26182_9_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_74 = T_26182_10_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_74 = T_26182_11_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_74 = T_26182_12_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_74 = T_26182_13_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_74 = T_26182_14_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_74 = T_26182_15_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_74 = T_26182_16_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_74 = T_26182_17_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_74 = T_26182_18_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_74 = T_26182_19_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_74 = T_26182_20_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_74 = T_26182_21_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_74 = T_26182_22_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_74 = T_26182_23_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_74 = T_26182_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_75 = T_26182_1_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_75 = T_26182_2_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_75 = T_26182_3_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_75 = T_26182_4_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_75 = T_26182_5_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_75 = T_26182_6_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_75 = T_26182_7_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_75 = T_26182_8_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_75 = T_26182_9_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_75 = T_26182_10_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_75 = T_26182_11_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_75 = T_26182_12_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_75 = T_26182_13_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_75 = T_26182_14_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_75 = T_26182_15_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_75 = T_26182_16_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_75 = T_26182_17_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_75 = T_26182_18_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_75 = T_26182_19_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_75 = T_26182_20_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_75 = T_26182_21_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_75 = T_26182_22_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_75 = T_26182_23_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_75 = T_26182_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_76 = T_26182_1_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_76 = T_26182_2_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_76 = T_26182_3_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_76 = T_26182_4_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_76 = T_26182_5_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_76 = T_26182_6_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_76 = T_26182_7_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_76 = T_26182_8_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_76 = T_26182_9_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_76 = T_26182_10_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_76 = T_26182_11_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_76 = T_26182_12_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_76 = T_26182_13_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_76 = T_26182_14_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_76 = T_26182_15_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_76 = T_26182_16_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_76 = T_26182_17_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_76 = T_26182_18_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_76 = T_26182_19_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_76 = T_26182_20_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_76 = T_26182_21_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_76 = T_26182_22_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_76 = T_26182_23_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_76 = T_26182_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_77 = T_26182_1_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_77 = T_26182_2_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_77 = T_26182_3_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_77 = T_26182_4_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_77 = T_26182_5_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_77 = T_26182_6_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_77 = T_26182_7_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_77 = T_26182_8_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_77 = T_26182_9_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_77 = T_26182_10_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_77 = T_26182_11_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_77 = T_26182_12_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_77 = T_26182_13_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_77 = T_26182_14_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_77 = T_26182_15_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_77 = T_26182_16_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_77 = T_26182_17_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_77 = T_26182_18_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_77 = T_26182_19_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_77 = T_26182_20_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_77 = T_26182_21_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_77 = T_26182_22_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_77 = T_26182_23_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_77 = T_26182_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_78 = T_26182_1_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_78 = T_26182_2_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_78 = T_26182_3_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_78 = T_26182_4_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_78 = T_26182_5_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_78 = T_26182_6_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_78 = T_26182_7_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_78 = T_26182_8_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_78 = T_26182_9_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_78 = T_26182_10_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_78 = T_26182_11_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_78 = T_26182_12_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_78 = T_26182_13_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_78 = T_26182_14_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_78 = T_26182_15_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_78 = T_26182_16_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_78 = T_26182_17_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_78 = T_26182_18_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_78 = T_26182_19_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_78 = T_26182_20_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_78 = T_26182_21_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_78 = T_26182_22_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_78 = T_26182_23_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_78 = T_26182_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_79 = T_26182_1_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_79 = T_26182_2_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_79 = T_26182_3_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_79 = T_26182_4_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_79 = T_26182_5_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_79 = T_26182_6_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_79 = T_26182_7_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_79 = T_26182_8_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_79 = T_26182_9_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_79 = T_26182_10_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_79 = T_26182_11_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_79 = T_26182_12_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_79 = T_26182_13_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_79 = T_26182_14_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_79 = T_26182_15_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_79 = T_26182_16_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_79 = T_26182_17_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_79 = T_26182_18_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_79 = T_26182_19_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_79 = T_26182_20_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_79 = T_26182_21_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_79 = T_26182_22_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_79 = T_26182_23_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_79 = T_26182_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_80 = T_26182_1_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_80 = T_26182_2_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_80 = T_26182_3_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_80 = T_26182_4_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_80 = T_26182_5_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_80 = T_26182_6_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_80 = T_26182_7_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_80 = T_26182_8_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_80 = T_26182_9_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_80 = T_26182_10_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_80 = T_26182_11_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_80 = T_26182_12_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_80 = T_26182_13_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_80 = T_26182_14_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_80 = T_26182_15_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_80 = T_26182_16_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_80 = T_26182_17_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_80 = T_26182_18_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_80 = T_26182_19_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_80 = T_26182_20_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_80 = T_26182_21_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_80 = T_26182_22_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_80 = T_26182_23_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_80 = T_26182_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_81 = T_26182_1_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_81 = T_26182_2_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_81 = T_26182_3_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_81 = T_26182_4_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_81 = T_26182_5_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_81 = T_26182_6_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_81 = T_26182_7_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_81 = T_26182_8_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_81 = T_26182_9_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_81 = T_26182_10_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_81 = T_26182_11_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_81 = T_26182_12_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_81 = T_26182_13_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_81 = T_26182_14_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_81 = T_26182_15_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_81 = T_26182_16_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_81 = T_26182_17_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_81 = T_26182_18_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_81 = T_26182_19_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_81 = T_26182_20_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_81 = T_26182_21_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_81 = T_26182_22_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_81 = T_26182_23_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_81 = T_26182_0_is_store;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_82 = T_26182_1_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_82 = T_26182_2_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_82 = T_26182_3_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_82 = T_26182_4_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_82 = T_26182_5_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_82 = T_26182_6_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_82 = T_26182_7_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_82 = T_26182_8_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_82 = T_26182_9_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_82 = T_26182_10_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_82 = T_26182_11_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_82 = T_26182_12_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_82 = T_26182_13_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_82 = T_26182_14_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_82 = T_26182_15_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_82 = T_26182_16_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_82 = T_26182_17_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_82 = T_26182_18_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_82 = T_26182_19_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_82 = T_26182_20_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_82 = T_26182_21_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_82 = T_26182_22_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_82 = T_26182_23_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_82 = T_26182_0_is_load;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_83 = T_26182_1_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_83 = T_26182_2_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_83 = T_26182_3_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_83 = T_26182_4_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_83 = T_26182_5_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_83 = T_26182_6_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_83 = T_26182_7_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_83 = T_26182_8_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_83 = T_26182_9_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_83 = T_26182_10_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_83 = T_26182_11_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_83 = T_26182_12_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_83 = T_26182_13_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_83 = T_26182_14_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_83 = T_26182_15_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_83 = T_26182_16_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_83 = T_26182_17_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_83 = T_26182_18_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_83 = T_26182_19_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_83 = T_26182_20_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_83 = T_26182_21_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_83 = T_26182_22_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_83 = T_26182_23_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_83 = T_26182_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  wire [5:0] _T_31993 = _io_get_pc_rob_idx_5to1 == 5'h17 ? 6'h0 : {1'h0, _io_get_pc_rob_idx_5to1} + 6'h1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:347:34, :967:16, util.scala:75:28, :76:{13,35}
  assign _T_1 = _T_31993 == 6'h17 ? T_23706_23 : _T_31993 == 6'h16 ? T_23706_22 : _T_31993 == 6'h15 ?
                T_23706_21 : _T_31993 == 6'h14 ? T_23706_20 : _T_31993 == 6'h13 ? T_23706_19 : _T_31993 ==
                6'h12 ? T_23706_18 : _T_31993 == 6'h11 ? T_23706_17 : _T_31993 == 6'h10 ? T_23706_16 :
                _T_31993 == 6'hF ? T_23706_15 : _T_31993 == 6'hE ? T_23706_14 : _T_31993 == 6'hD ?
                T_23706_13 : _T_31993 == 6'hC ? T_23706_12 : _T_31993 == 6'hB ? T_23706_11 : _T_31993 ==
                6'hA ? T_23706_10 : _T_31993 == 6'h9 ? T_23706_9 : _T_31993 == 6'h8 ? T_23706_8 : _T_31993
                == 6'h7 ? T_23706_7 : _T_31993 == 6'h6 ? T_23706_6 : _T_31993 == 6'h5 ? T_23706_5 :
                _T_31993 == 6'h4 ? T_23706_4 : _T_31993 == 6'h3 ? T_23706_3 : _T_31993 == 6'h2 ? T_23706_2
                : _T_31993 == 6'h1 ? T_23706_1 : T_23706_0;	// rob.scala:347:34, :509:28, :967:16
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_84 = T_23706_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_84 = T_23706_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_84 = T_23706_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_84 = T_23706_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_84 = T_23706_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_84 = T_23706_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_84 = T_23706_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_84 = T_23706_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_84 = T_23706_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_84 = T_23706_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_84 = T_23706_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_84 = T_23706_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_84 = T_23706_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_84 = T_23706_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_84 = T_23706_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_84 = T_23706_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_84 = T_23706_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_84 = T_23706_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_84 = T_23706_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_84 = T_23706_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_84 = T_23706_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_84 = T_23706_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_84 = T_23706_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_84 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_85 = T_26182_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_85 = T_26182_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_85 = T_26182_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_85 = T_26182_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_85 = T_26182_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_85 = T_26182_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_85 = T_26182_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_85 = T_26182_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_85 = T_26182_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_85 = T_26182_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_85 = T_26182_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_85 = T_26182_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_85 = T_26182_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_85 = T_26182_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_85 = T_26182_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_85 = T_26182_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_85 = T_26182_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_85 = T_26182_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_85 = T_26182_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_85 = T_26182_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_85 = T_26182_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_85 = T_26182_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_85 = T_26182_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_85 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_86 = T_26182_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_86 = T_26182_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_86 = T_26182_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_86 = T_26182_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_86 = T_26182_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_86 = T_26182_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_86 = T_26182_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_86 = T_26182_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_86 = T_26182_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_86 = T_26182_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_86 = T_26182_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_86 = T_26182_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_86 = T_26182_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_86 = T_26182_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_86 = T_26182_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_86 = T_26182_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_86 = T_26182_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_86 = T_26182_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_86 = T_26182_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_86 = T_26182_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_86 = T_26182_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_86 = T_26182_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_86 = T_26182_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_86 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_87 = T_23706_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_87 = T_23706_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_87 = T_23706_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_87 = T_23706_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_87 = T_23706_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_87 = T_23706_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_87 = T_23706_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_87 = T_23706_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_87 = T_23706_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_87 = T_23706_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_87 = T_23706_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_87 = T_23706_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_87 = T_23706_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_87 = T_23706_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_87 = T_23706_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_87 = T_23706_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_87 = T_23706_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_87 = T_23706_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_87 = T_23706_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_87 = T_23706_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_87 = T_23706_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_87 = T_23706_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_87 = T_23706_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_87 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_88 = T_26182_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_88 = T_26182_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_88 = T_26182_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_88 = T_26182_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_88 = T_26182_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_88 = T_26182_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_88 = T_26182_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_88 = T_26182_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_88 = T_26182_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_88 = T_26182_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_88 = T_26182_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_88 = T_26182_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_88 = T_26182_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_88 = T_26182_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_88 = T_26182_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_88 = T_26182_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_88 = T_26182_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_88 = T_26182_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_88 = T_26182_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_88 = T_26182_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_88 = T_26182_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_88 = T_26182_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_88 = T_26182_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_88 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_89 = T_26182_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_89 = T_26182_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_89 = T_26182_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_89 = T_26182_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_89 = T_26182_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_89 = T_26182_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_89 = T_26182_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_89 = T_26182_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_89 = T_26182_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_89 = T_26182_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_89 = T_26182_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_89 = T_26182_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_89 = T_26182_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_89 = T_26182_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_89 = T_26182_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_89 = T_26182_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_89 = T_26182_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_89 = T_26182_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_89 = T_26182_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_89 = T_26182_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_89 = T_26182_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_89 = T_26182_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_89 = T_26182_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_89 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_90 = T_23706_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_90 = T_23706_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_90 = T_23706_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_90 = T_23706_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_90 = T_23706_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_90 = T_23706_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_90 = T_23706_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_90 = T_23706_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_90 = T_23706_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_90 = T_23706_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_90 = T_23706_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_90 = T_23706_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_90 = T_23706_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_90 = T_23706_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_90 = T_23706_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_90 = T_23706_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_90 = T_23706_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_90 = T_23706_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_90 = T_23706_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_90 = T_23706_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_90 = T_23706_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_90 = T_23706_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_90 = T_23706_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_90 = T_23706_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_91 = T_26182_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_91 = T_26182_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_91 = T_26182_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_91 = T_26182_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_91 = T_26182_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_91 = T_26182_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_91 = T_26182_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_91 = T_26182_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_91 = T_26182_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_91 = T_26182_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_91 = T_26182_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_91 = T_26182_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_91 = T_26182_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_91 = T_26182_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_91 = T_26182_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_91 = T_26182_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_91 = T_26182_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_91 = T_26182_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_91 = T_26182_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_91 = T_26182_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_91 = T_26182_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_91 = T_26182_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_91 = T_26182_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_91 = T_26182_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_92 = T_26182_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_92 = T_26182_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_92 = T_26182_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_92 = T_26182_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_92 = T_26182_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_92 = T_26182_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_92 = T_26182_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_92 = T_26182_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_92 = T_26182_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_92 = T_26182_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_92 = T_26182_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_92 = T_26182_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_92 = T_26182_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_92 = T_26182_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_92 = T_26182_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_92 = T_26182_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_92 = T_26182_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_92 = T_26182_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_92 = T_26182_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_92 = T_26182_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_92 = T_26182_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_92 = T_26182_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_92 = T_26182_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_92 = T_26182_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:347:34, :355:47
    casez (rob_tail)	// rob.scala:192:32, :347:34, :355:47
      5'b00000:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b00001:
        casez_tmp_93 = T_35634_1;	// rob.scala:347:34, :355:47
      5'b00010:
        casez_tmp_93 = T_35634_2;	// rob.scala:347:34, :355:47
      5'b00011:
        casez_tmp_93 = T_35634_3;	// rob.scala:347:34, :355:47
      5'b00100:
        casez_tmp_93 = T_35634_4;	// rob.scala:347:34, :355:47
      5'b00101:
        casez_tmp_93 = T_35634_5;	// rob.scala:347:34, :355:47
      5'b00110:
        casez_tmp_93 = T_35634_6;	// rob.scala:347:34, :355:47
      5'b00111:
        casez_tmp_93 = T_35634_7;	// rob.scala:347:34, :355:47
      5'b01000:
        casez_tmp_93 = T_35634_8;	// rob.scala:347:34, :355:47
      5'b01001:
        casez_tmp_93 = T_35634_9;	// rob.scala:347:34, :355:47
      5'b01010:
        casez_tmp_93 = T_35634_10;	// rob.scala:347:34, :355:47
      5'b01011:
        casez_tmp_93 = T_35634_11;	// rob.scala:347:34, :355:47
      5'b01100:
        casez_tmp_93 = T_35634_12;	// rob.scala:347:34, :355:47
      5'b01101:
        casez_tmp_93 = T_35634_13;	// rob.scala:347:34, :355:47
      5'b01110:
        casez_tmp_93 = T_35634_14;	// rob.scala:347:34, :355:47
      5'b01111:
        casez_tmp_93 = T_35634_15;	// rob.scala:347:34, :355:47
      5'b10000:
        casez_tmp_93 = T_35634_16;	// rob.scala:347:34, :355:47
      5'b10001:
        casez_tmp_93 = T_35634_17;	// rob.scala:347:34, :355:47
      5'b10010:
        casez_tmp_93 = T_35634_18;	// rob.scala:347:34, :355:47
      5'b10011:
        casez_tmp_93 = T_35634_19;	// rob.scala:347:34, :355:47
      5'b10100:
        casez_tmp_93 = T_35634_20;	// rob.scala:347:34, :355:47
      5'b10101:
        casez_tmp_93 = T_35634_21;	// rob.scala:347:34, :355:47
      5'b10110:
        casez_tmp_93 = T_35634_22;	// rob.scala:347:34, :355:47
      5'b10111:
        casez_tmp_93 = T_35634_23;	// rob.scala:347:34, :355:47
      5'b11000:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11001:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11010:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11011:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11100:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11101:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      5'b11110:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
      default:
        casez_tmp_93 = T_35634_0;	// rob.scala:347:34, :355:47
    endcase	// rob.scala:192:32, :347:34, :355:47
  end // always @(*)
  always @(*) begin	// rob.scala:433:51
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51
      5'b00000:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b00001:
        casez_tmp_94 = T_35634_1;	// rob.scala:347:34, :433:51
      5'b00010:
        casez_tmp_94 = T_35634_2;	// rob.scala:347:34, :433:51
      5'b00011:
        casez_tmp_94 = T_35634_3;	// rob.scala:347:34, :433:51
      5'b00100:
        casez_tmp_94 = T_35634_4;	// rob.scala:347:34, :433:51
      5'b00101:
        casez_tmp_94 = T_35634_5;	// rob.scala:347:34, :433:51
      5'b00110:
        casez_tmp_94 = T_35634_6;	// rob.scala:347:34, :433:51
      5'b00111:
        casez_tmp_94 = T_35634_7;	// rob.scala:347:34, :433:51
      5'b01000:
        casez_tmp_94 = T_35634_8;	// rob.scala:347:34, :433:51
      5'b01001:
        casez_tmp_94 = T_35634_9;	// rob.scala:347:34, :433:51
      5'b01010:
        casez_tmp_94 = T_35634_10;	// rob.scala:347:34, :433:51
      5'b01011:
        casez_tmp_94 = T_35634_11;	// rob.scala:347:34, :433:51
      5'b01100:
        casez_tmp_94 = T_35634_12;	// rob.scala:347:34, :433:51
      5'b01101:
        casez_tmp_94 = T_35634_13;	// rob.scala:347:34, :433:51
      5'b01110:
        casez_tmp_94 = T_35634_14;	// rob.scala:347:34, :433:51
      5'b01111:
        casez_tmp_94 = T_35634_15;	// rob.scala:347:34, :433:51
      5'b10000:
        casez_tmp_94 = T_35634_16;	// rob.scala:347:34, :433:51
      5'b10001:
        casez_tmp_94 = T_35634_17;	// rob.scala:347:34, :433:51
      5'b10010:
        casez_tmp_94 = T_35634_18;	// rob.scala:347:34, :433:51
      5'b10011:
        casez_tmp_94 = T_35634_19;	// rob.scala:347:34, :433:51
      5'b10100:
        casez_tmp_94 = T_35634_20;	// rob.scala:347:34, :433:51
      5'b10101:
        casez_tmp_94 = T_35634_21;	// rob.scala:347:34, :433:51
      5'b10110:
        casez_tmp_94 = T_35634_22;	// rob.scala:347:34, :433:51
      5'b10111:
        casez_tmp_94 = T_35634_23;	// rob.scala:347:34, :433:51
      5'b11000:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11001:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11010:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11011:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11100:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11101:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      5'b11110:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
      default:
        casez_tmp_94 = T_35634_0;	// rob.scala:347:34, :433:51
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51
  end // always @(*)
  wire _T_41018 = casez_tmp_94 & T_40239_R0_data;	// rob.scala:339:30, :433:51
  always @(*) begin	// rob.scala:451:58
    casez (_T_2)	// rob.scala:451:58
      5'b00000:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b00001:
        casez_tmp_95 = T_35634_1;	// rob.scala:347:34, :451:58
      5'b00010:
        casez_tmp_95 = T_35634_2;	// rob.scala:347:34, :451:58
      5'b00011:
        casez_tmp_95 = T_35634_3;	// rob.scala:347:34, :451:58
      5'b00100:
        casez_tmp_95 = T_35634_4;	// rob.scala:347:34, :451:58
      5'b00101:
        casez_tmp_95 = T_35634_5;	// rob.scala:347:34, :451:58
      5'b00110:
        casez_tmp_95 = T_35634_6;	// rob.scala:347:34, :451:58
      5'b00111:
        casez_tmp_95 = T_35634_7;	// rob.scala:347:34, :451:58
      5'b01000:
        casez_tmp_95 = T_35634_8;	// rob.scala:347:34, :451:58
      5'b01001:
        casez_tmp_95 = T_35634_9;	// rob.scala:347:34, :451:58
      5'b01010:
        casez_tmp_95 = T_35634_10;	// rob.scala:347:34, :451:58
      5'b01011:
        casez_tmp_95 = T_35634_11;	// rob.scala:347:34, :451:58
      5'b01100:
        casez_tmp_95 = T_35634_12;	// rob.scala:347:34, :451:58
      5'b01101:
        casez_tmp_95 = T_35634_13;	// rob.scala:347:34, :451:58
      5'b01110:
        casez_tmp_95 = T_35634_14;	// rob.scala:347:34, :451:58
      5'b01111:
        casez_tmp_95 = T_35634_15;	// rob.scala:347:34, :451:58
      5'b10000:
        casez_tmp_95 = T_35634_16;	// rob.scala:347:34, :451:58
      5'b10001:
        casez_tmp_95 = T_35634_17;	// rob.scala:347:34, :451:58
      5'b10010:
        casez_tmp_95 = T_35634_18;	// rob.scala:347:34, :451:58
      5'b10011:
        casez_tmp_95 = T_35634_19;	// rob.scala:347:34, :451:58
      5'b10100:
        casez_tmp_95 = T_35634_20;	// rob.scala:347:34, :451:58
      5'b10101:
        casez_tmp_95 = T_35634_21;	// rob.scala:347:34, :451:58
      5'b10110:
        casez_tmp_95 = T_35634_22;	// rob.scala:347:34, :451:58
      5'b10111:
        casez_tmp_95 = T_35634_23;	// rob.scala:347:34, :451:58
      5'b11000:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11001:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11010:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11011:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11100:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11101:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      5'b11110:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
      default:
        casez_tmp_95 = T_35634_0;	// rob.scala:347:34, :451:58
    endcase	// rob.scala:451:58
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_96 = T_38110_1_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_96 = T_38110_2_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_96 = T_38110_3_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_96 = T_38110_4_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_96 = T_38110_5_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_96 = T_38110_6_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_96 = T_38110_7_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_96 = T_38110_8_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_96 = T_38110_9_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_96 = T_38110_10_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_96 = T_38110_11_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_96 = T_38110_12_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_96 = T_38110_13_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_96 = T_38110_14_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_96 = T_38110_15_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_96 = T_38110_16_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_96 = T_38110_17_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_96 = T_38110_18_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_96 = T_38110_19_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_96 = T_38110_20_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_96 = T_38110_21_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_96 = T_38110_22_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_96 = T_38110_23_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_96 = T_38110_0_valid;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_97 = T_38110_1_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_97 = T_38110_2_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_97 = T_38110_3_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_97 = T_38110_4_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_97 = T_38110_5_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_97 = T_38110_6_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_97 = T_38110_7_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_97 = T_38110_8_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_97 = T_38110_9_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_97 = T_38110_10_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_97 = T_38110_11_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_97 = T_38110_12_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_97 = T_38110_13_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_97 = T_38110_14_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_97 = T_38110_15_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_97 = T_38110_16_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_97 = T_38110_17_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_97 = T_38110_18_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_97 = T_38110_19_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_97 = T_38110_20_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_97 = T_38110_21_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_97 = T_38110_22_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_97 = T_38110_23_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_97 = T_38110_0_iw_state;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_98 = T_38110_1_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_98 = T_38110_2_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_98 = T_38110_3_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_98 = T_38110_4_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_98 = T_38110_5_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_98 = T_38110_6_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_98 = T_38110_7_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_98 = T_38110_8_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_98 = T_38110_9_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_98 = T_38110_10_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_98 = T_38110_11_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_98 = T_38110_12_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_98 = T_38110_13_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_98 = T_38110_14_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_98 = T_38110_15_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_98 = T_38110_16_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_98 = T_38110_17_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_98 = T_38110_18_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_98 = T_38110_19_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_98 = T_38110_20_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_98 = T_38110_21_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_98 = T_38110_22_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_98 = T_38110_23_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_98 = T_38110_0_uopc;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_99 = T_38110_1_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_99 = T_38110_2_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_99 = T_38110_3_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_99 = T_38110_4_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_99 = T_38110_5_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_99 = T_38110_6_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_99 = T_38110_7_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_99 = T_38110_8_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_99 = T_38110_9_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_99 = T_38110_10_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_99 = T_38110_11_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_99 = T_38110_12_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_99 = T_38110_13_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_99 = T_38110_14_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_99 = T_38110_15_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_99 = T_38110_16_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_99 = T_38110_17_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_99 = T_38110_18_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_99 = T_38110_19_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_99 = T_38110_20_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_99 = T_38110_21_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_99 = T_38110_22_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_99 = T_38110_23_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_99 = T_38110_0_inst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_100 = T_38110_1_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_100 = T_38110_2_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_100 = T_38110_3_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_100 = T_38110_4_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_100 = T_38110_5_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_100 = T_38110_6_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_100 = T_38110_7_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_100 = T_38110_8_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_100 = T_38110_9_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_100 = T_38110_10_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_100 = T_38110_11_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_100 = T_38110_12_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_100 = T_38110_13_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_100 = T_38110_14_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_100 = T_38110_15_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_100 = T_38110_16_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_100 = T_38110_17_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_100 = T_38110_18_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_100 = T_38110_19_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_100 = T_38110_20_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_100 = T_38110_21_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_100 = T_38110_22_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_100 = T_38110_23_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_100 = T_38110_0_pc;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_101 = T_38110_1_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_101 = T_38110_2_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_101 = T_38110_3_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_101 = T_38110_4_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_101 = T_38110_5_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_101 = T_38110_6_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_101 = T_38110_7_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_101 = T_38110_8_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_101 = T_38110_9_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_101 = T_38110_10_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_101 = T_38110_11_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_101 = T_38110_12_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_101 = T_38110_13_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_101 = T_38110_14_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_101 = T_38110_15_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_101 = T_38110_16_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_101 = T_38110_17_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_101 = T_38110_18_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_101 = T_38110_19_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_101 = T_38110_20_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_101 = T_38110_21_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_101 = T_38110_22_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_101 = T_38110_23_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_101 = T_38110_0_fu_code;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_102 = T_38110_1_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_102 = T_38110_2_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_102 = T_38110_3_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_102 = T_38110_4_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_102 = T_38110_5_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_102 = T_38110_6_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_102 = T_38110_7_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_102 = T_38110_8_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_102 = T_38110_9_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_102 = T_38110_10_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_102 = T_38110_11_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_102 = T_38110_12_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_102 = T_38110_13_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_102 = T_38110_14_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_102 = T_38110_15_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_102 = T_38110_16_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_102 = T_38110_17_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_102 = T_38110_18_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_102 = T_38110_19_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_102 = T_38110_20_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_102 = T_38110_21_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_102 = T_38110_22_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_102 = T_38110_23_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_102 = T_38110_0_ctrl_br_type;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_103 = T_38110_1_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_103 = T_38110_2_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_103 = T_38110_3_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_103 = T_38110_4_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_103 = T_38110_5_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_103 = T_38110_6_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_103 = T_38110_7_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_103 = T_38110_8_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_103 = T_38110_9_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_103 = T_38110_10_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_103 = T_38110_11_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_103 = T_38110_12_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_103 = T_38110_13_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_103 = T_38110_14_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_103 = T_38110_15_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_103 = T_38110_16_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_103 = T_38110_17_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_103 = T_38110_18_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_103 = T_38110_19_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_103 = T_38110_20_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_103 = T_38110_21_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_103 = T_38110_22_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_103 = T_38110_23_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_103 = T_38110_0_ctrl_op1_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_104 = T_38110_1_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_104 = T_38110_2_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_104 = T_38110_3_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_104 = T_38110_4_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_104 = T_38110_5_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_104 = T_38110_6_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_104 = T_38110_7_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_104 = T_38110_8_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_104 = T_38110_9_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_104 = T_38110_10_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_104 = T_38110_11_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_104 = T_38110_12_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_104 = T_38110_13_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_104 = T_38110_14_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_104 = T_38110_15_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_104 = T_38110_16_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_104 = T_38110_17_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_104 = T_38110_18_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_104 = T_38110_19_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_104 = T_38110_20_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_104 = T_38110_21_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_104 = T_38110_22_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_104 = T_38110_23_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_104 = T_38110_0_ctrl_op2_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_105 = T_38110_1_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_105 = T_38110_2_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_105 = T_38110_3_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_105 = T_38110_4_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_105 = T_38110_5_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_105 = T_38110_6_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_105 = T_38110_7_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_105 = T_38110_8_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_105 = T_38110_9_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_105 = T_38110_10_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_105 = T_38110_11_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_105 = T_38110_12_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_105 = T_38110_13_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_105 = T_38110_14_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_105 = T_38110_15_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_105 = T_38110_16_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_105 = T_38110_17_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_105 = T_38110_18_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_105 = T_38110_19_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_105 = T_38110_20_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_105 = T_38110_21_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_105 = T_38110_22_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_105 = T_38110_23_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_105 = T_38110_0_ctrl_imm_sel;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_106 = T_38110_1_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_106 = T_38110_2_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_106 = T_38110_3_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_106 = T_38110_4_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_106 = T_38110_5_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_106 = T_38110_6_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_106 = T_38110_7_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_106 = T_38110_8_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_106 = T_38110_9_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_106 = T_38110_10_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_106 = T_38110_11_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_106 = T_38110_12_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_106 = T_38110_13_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_106 = T_38110_14_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_106 = T_38110_15_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_106 = T_38110_16_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_106 = T_38110_17_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_106 = T_38110_18_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_106 = T_38110_19_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_106 = T_38110_20_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_106 = T_38110_21_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_106 = T_38110_22_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_106 = T_38110_23_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_106 = T_38110_0_ctrl_op_fcn;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_107 = T_38110_1_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_107 = T_38110_2_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_107 = T_38110_3_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_107 = T_38110_4_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_107 = T_38110_5_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_107 = T_38110_6_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_107 = T_38110_7_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_107 = T_38110_8_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_107 = T_38110_9_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_107 = T_38110_10_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_107 = T_38110_11_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_107 = T_38110_12_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_107 = T_38110_13_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_107 = T_38110_14_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_107 = T_38110_15_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_107 = T_38110_16_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_107 = T_38110_17_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_107 = T_38110_18_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_107 = T_38110_19_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_107 = T_38110_20_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_107 = T_38110_21_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_107 = T_38110_22_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_107 = T_38110_23_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_107 = T_38110_0_ctrl_fcn_dw;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_108 = T_38110_1_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_108 = T_38110_2_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_108 = T_38110_3_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_108 = T_38110_4_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_108 = T_38110_5_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_108 = T_38110_6_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_108 = T_38110_7_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_108 = T_38110_8_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_108 = T_38110_9_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_108 = T_38110_10_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_108 = T_38110_11_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_108 = T_38110_12_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_108 = T_38110_13_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_108 = T_38110_14_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_108 = T_38110_15_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_108 = T_38110_16_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_108 = T_38110_17_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_108 = T_38110_18_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_108 = T_38110_19_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_108 = T_38110_20_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_108 = T_38110_21_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_108 = T_38110_22_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_108 = T_38110_23_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_108 = T_38110_0_ctrl_rf_wen;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_109 = T_38110_1_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_109 = T_38110_2_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_109 = T_38110_3_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_109 = T_38110_4_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_109 = T_38110_5_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_109 = T_38110_6_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_109 = T_38110_7_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_109 = T_38110_8_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_109 = T_38110_9_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_109 = T_38110_10_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_109 = T_38110_11_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_109 = T_38110_12_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_109 = T_38110_13_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_109 = T_38110_14_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_109 = T_38110_15_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_109 = T_38110_16_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_109 = T_38110_17_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_109 = T_38110_18_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_109 = T_38110_19_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_109 = T_38110_20_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_109 = T_38110_21_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_109 = T_38110_22_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_109 = T_38110_23_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_109 = T_38110_0_ctrl_csr_cmd;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_110 = T_38110_1_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_110 = T_38110_2_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_110 = T_38110_3_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_110 = T_38110_4_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_110 = T_38110_5_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_110 = T_38110_6_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_110 = T_38110_7_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_110 = T_38110_8_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_110 = T_38110_9_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_110 = T_38110_10_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_110 = T_38110_11_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_110 = T_38110_12_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_110 = T_38110_13_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_110 = T_38110_14_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_110 = T_38110_15_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_110 = T_38110_16_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_110 = T_38110_17_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_110 = T_38110_18_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_110 = T_38110_19_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_110 = T_38110_20_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_110 = T_38110_21_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_110 = T_38110_22_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_110 = T_38110_23_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_110 = T_38110_0_ctrl_is_load;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_111 = T_38110_1_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_111 = T_38110_2_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_111 = T_38110_3_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_111 = T_38110_4_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_111 = T_38110_5_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_111 = T_38110_6_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_111 = T_38110_7_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_111 = T_38110_8_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_111 = T_38110_9_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_111 = T_38110_10_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_111 = T_38110_11_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_111 = T_38110_12_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_111 = T_38110_13_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_111 = T_38110_14_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_111 = T_38110_15_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_111 = T_38110_16_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_111 = T_38110_17_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_111 = T_38110_18_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_111 = T_38110_19_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_111 = T_38110_20_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_111 = T_38110_21_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_111 = T_38110_22_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_111 = T_38110_23_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_111 = T_38110_0_ctrl_is_sta;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_112 = T_38110_1_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_112 = T_38110_2_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_112 = T_38110_3_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_112 = T_38110_4_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_112 = T_38110_5_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_112 = T_38110_6_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_112 = T_38110_7_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_112 = T_38110_8_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_112 = T_38110_9_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_112 = T_38110_10_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_112 = T_38110_11_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_112 = T_38110_12_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_112 = T_38110_13_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_112 = T_38110_14_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_112 = T_38110_15_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_112 = T_38110_16_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_112 = T_38110_17_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_112 = T_38110_18_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_112 = T_38110_19_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_112 = T_38110_20_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_112 = T_38110_21_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_112 = T_38110_22_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_112 = T_38110_23_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_112 = T_38110_0_ctrl_is_std;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_113 = T_38110_1_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_113 = T_38110_2_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_113 = T_38110_3_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_113 = T_38110_4_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_113 = T_38110_5_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_113 = T_38110_6_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_113 = T_38110_7_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_113 = T_38110_8_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_113 = T_38110_9_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_113 = T_38110_10_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_113 = T_38110_11_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_113 = T_38110_12_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_113 = T_38110_13_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_113 = T_38110_14_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_113 = T_38110_15_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_113 = T_38110_16_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_113 = T_38110_17_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_113 = T_38110_18_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_113 = T_38110_19_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_113 = T_38110_20_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_113 = T_38110_21_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_113 = T_38110_22_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_113 = T_38110_23_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_113 = T_38110_0_wakeup_delay;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_114 = T_38110_1_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_114 = T_38110_2_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_114 = T_38110_3_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_114 = T_38110_4_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_114 = T_38110_5_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_114 = T_38110_6_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_114 = T_38110_7_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_114 = T_38110_8_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_114 = T_38110_9_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_114 = T_38110_10_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_114 = T_38110_11_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_114 = T_38110_12_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_114 = T_38110_13_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_114 = T_38110_14_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_114 = T_38110_15_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_114 = T_38110_16_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_114 = T_38110_17_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_114 = T_38110_18_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_114 = T_38110_19_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_114 = T_38110_20_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_114 = T_38110_21_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_114 = T_38110_22_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_114 = T_38110_23_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_114 = T_38110_0_allocate_brtag;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_115 = T_38110_1_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_115 = T_38110_2_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_115 = T_38110_3_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_115 = T_38110_4_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_115 = T_38110_5_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_115 = T_38110_6_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_115 = T_38110_7_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_115 = T_38110_8_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_115 = T_38110_9_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_115 = T_38110_10_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_115 = T_38110_11_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_115 = T_38110_12_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_115 = T_38110_13_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_115 = T_38110_14_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_115 = T_38110_15_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_115 = T_38110_16_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_115 = T_38110_17_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_115 = T_38110_18_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_115 = T_38110_19_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_115 = T_38110_20_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_115 = T_38110_21_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_115 = T_38110_22_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_115 = T_38110_23_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_115 = T_38110_0_is_br_or_jmp;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_116 = T_38110_1_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_116 = T_38110_2_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_116 = T_38110_3_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_116 = T_38110_4_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_116 = T_38110_5_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_116 = T_38110_6_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_116 = T_38110_7_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_116 = T_38110_8_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_116 = T_38110_9_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_116 = T_38110_10_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_116 = T_38110_11_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_116 = T_38110_12_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_116 = T_38110_13_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_116 = T_38110_14_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_116 = T_38110_15_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_116 = T_38110_16_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_116 = T_38110_17_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_116 = T_38110_18_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_116 = T_38110_19_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_116 = T_38110_20_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_116 = T_38110_21_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_116 = T_38110_22_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_116 = T_38110_23_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_116 = T_38110_0_is_jump;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_117 = T_38110_1_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_117 = T_38110_2_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_117 = T_38110_3_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_117 = T_38110_4_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_117 = T_38110_5_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_117 = T_38110_6_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_117 = T_38110_7_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_117 = T_38110_8_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_117 = T_38110_9_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_117 = T_38110_10_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_117 = T_38110_11_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_117 = T_38110_12_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_117 = T_38110_13_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_117 = T_38110_14_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_117 = T_38110_15_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_117 = T_38110_16_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_117 = T_38110_17_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_117 = T_38110_18_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_117 = T_38110_19_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_117 = T_38110_20_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_117 = T_38110_21_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_117 = T_38110_22_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_117 = T_38110_23_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_117 = T_38110_0_is_jal;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_118 = T_38110_1_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_118 = T_38110_2_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_118 = T_38110_3_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_118 = T_38110_4_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_118 = T_38110_5_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_118 = T_38110_6_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_118 = T_38110_7_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_118 = T_38110_8_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_118 = T_38110_9_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_118 = T_38110_10_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_118 = T_38110_11_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_118 = T_38110_12_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_118 = T_38110_13_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_118 = T_38110_14_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_118 = T_38110_15_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_118 = T_38110_16_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_118 = T_38110_17_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_118 = T_38110_18_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_118 = T_38110_19_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_118 = T_38110_20_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_118 = T_38110_21_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_118 = T_38110_22_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_118 = T_38110_23_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_118 = T_38110_0_is_ret;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_119 = T_38110_1_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_119 = T_38110_2_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_119 = T_38110_3_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_119 = T_38110_4_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_119 = T_38110_5_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_119 = T_38110_6_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_119 = T_38110_7_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_119 = T_38110_8_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_119 = T_38110_9_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_119 = T_38110_10_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_119 = T_38110_11_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_119 = T_38110_12_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_119 = T_38110_13_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_119 = T_38110_14_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_119 = T_38110_15_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_119 = T_38110_16_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_119 = T_38110_17_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_119 = T_38110_18_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_119 = T_38110_19_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_119 = T_38110_20_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_119 = T_38110_21_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_119 = T_38110_22_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_119 = T_38110_23_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_119 = T_38110_0_is_call;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_120 = T_38110_1_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_120 = T_38110_2_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_120 = T_38110_3_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_120 = T_38110_4_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_120 = T_38110_5_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_120 = T_38110_6_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_120 = T_38110_7_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_120 = T_38110_8_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_120 = T_38110_9_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_120 = T_38110_10_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_120 = T_38110_11_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_120 = T_38110_12_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_120 = T_38110_13_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_120 = T_38110_14_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_120 = T_38110_15_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_120 = T_38110_16_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_120 = T_38110_17_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_120 = T_38110_18_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_120 = T_38110_19_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_120 = T_38110_20_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_120 = T_38110_21_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_120 = T_38110_22_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_120 = T_38110_23_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_120 = T_38110_0_br_mask;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_121 = T_38110_1_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_121 = T_38110_2_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_121 = T_38110_3_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_121 = T_38110_4_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_121 = T_38110_5_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_121 = T_38110_6_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_121 = T_38110_7_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_121 = T_38110_8_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_121 = T_38110_9_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_121 = T_38110_10_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_121 = T_38110_11_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_121 = T_38110_12_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_121 = T_38110_13_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_121 = T_38110_14_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_121 = T_38110_15_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_121 = T_38110_16_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_121 = T_38110_17_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_121 = T_38110_18_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_121 = T_38110_19_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_121 = T_38110_20_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_121 = T_38110_21_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_121 = T_38110_22_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_121 = T_38110_23_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_121 = T_38110_0_br_tag;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_122 = T_38110_1_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_122 = T_38110_2_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_122 = T_38110_3_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_122 = T_38110_4_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_122 = T_38110_5_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_122 = T_38110_6_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_122 = T_38110_7_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_122 = T_38110_8_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_122 = T_38110_9_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_122 = T_38110_10_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_122 = T_38110_11_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_122 = T_38110_12_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_122 = T_38110_13_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_122 = T_38110_14_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_122 = T_38110_15_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_122 = T_38110_16_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_122 = T_38110_17_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_122 = T_38110_18_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_122 = T_38110_19_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_122 = T_38110_20_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_122 = T_38110_21_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_122 = T_38110_22_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_122 = T_38110_23_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_122 = T_38110_0_br_prediction_bpd_predict_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_123 = T_38110_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_123 = T_38110_2_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_123 = T_38110_3_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_123 = T_38110_4_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_123 = T_38110_5_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_123 = T_38110_6_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_123 = T_38110_7_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_123 = T_38110_8_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_123 = T_38110_9_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_123 = T_38110_10_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_123 = T_38110_11_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_123 = T_38110_12_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_123 = T_38110_13_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_123 = T_38110_14_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_123 = T_38110_15_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_123 = T_38110_16_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_123 = T_38110_17_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_123 = T_38110_18_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_123 = T_38110_19_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_123 = T_38110_20_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_123 = T_38110_21_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_123 = T_38110_22_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_123 = T_38110_23_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_123 = T_38110_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_124 = T_38110_1_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_124 = T_38110_2_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_124 = T_38110_3_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_124 = T_38110_4_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_124 = T_38110_5_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_124 = T_38110_6_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_124 = T_38110_7_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_124 = T_38110_8_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_124 = T_38110_9_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_124 = T_38110_10_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_124 = T_38110_11_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_124 = T_38110_12_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_124 = T_38110_13_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_124 = T_38110_14_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_124 = T_38110_15_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_124 = T_38110_16_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_124 = T_38110_17_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_124 = T_38110_18_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_124 = T_38110_19_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_124 = T_38110_20_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_124 = T_38110_21_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_124 = T_38110_22_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_124 = T_38110_23_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_124 = T_38110_0_br_prediction_btb_hit;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_125 = T_38110_1_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_125 = T_38110_2_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_125 = T_38110_3_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_125 = T_38110_4_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_125 = T_38110_5_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_125 = T_38110_6_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_125 = T_38110_7_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_125 = T_38110_8_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_125 = T_38110_9_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_125 = T_38110_10_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_125 = T_38110_11_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_125 = T_38110_12_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_125 = T_38110_13_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_125 = T_38110_14_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_125 = T_38110_15_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_125 = T_38110_16_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_125 = T_38110_17_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_125 = T_38110_18_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_125 = T_38110_19_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_125 = T_38110_20_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_125 = T_38110_21_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_125 = T_38110_22_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_125 = T_38110_23_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_125 = T_38110_0_br_prediction_btb_predicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_126 = T_38110_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_126 = T_38110_2_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_126 = T_38110_3_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_126 = T_38110_4_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_126 = T_38110_5_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_126 = T_38110_6_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_126 = T_38110_7_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_126 = T_38110_8_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_126 = T_38110_9_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_126 = T_38110_10_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_126 = T_38110_11_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_126 = T_38110_12_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_126 = T_38110_13_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_126 = T_38110_14_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_126 = T_38110_15_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_126 = T_38110_16_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_126 = T_38110_17_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_126 = T_38110_18_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_126 = T_38110_19_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_126 = T_38110_20_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_126 = T_38110_21_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_126 = T_38110_22_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_126 = T_38110_23_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_126 = T_38110_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_127 = T_38110_1_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_127 = T_38110_2_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_127 = T_38110_3_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_127 = T_38110_4_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_127 = T_38110_5_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_127 = T_38110_6_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_127 = T_38110_7_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_127 = T_38110_8_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_127 = T_38110_9_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_127 = T_38110_10_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_127 = T_38110_11_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_127 = T_38110_12_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_127 = T_38110_13_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_127 = T_38110_14_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_127 = T_38110_15_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_127 = T_38110_16_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_127 = T_38110_17_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_127 = T_38110_18_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_127 = T_38110_19_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_127 = T_38110_20_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_127 = T_38110_21_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_127 = T_38110_22_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_127 = T_38110_23_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_127 = T_38110_0_stat_brjmp_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_128 = T_38110_1_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_128 = T_38110_2_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_128 = T_38110_3_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_128 = T_38110_4_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_128 = T_38110_5_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_128 = T_38110_6_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_128 = T_38110_7_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_128 = T_38110_8_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_128 = T_38110_9_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_128 = T_38110_10_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_128 = T_38110_11_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_128 = T_38110_12_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_128 = T_38110_13_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_128 = T_38110_14_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_128 = T_38110_15_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_128 = T_38110_16_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_128 = T_38110_17_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_128 = T_38110_18_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_128 = T_38110_19_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_128 = T_38110_20_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_128 = T_38110_21_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_128 = T_38110_22_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_128 = T_38110_23_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_128 = T_38110_0_stat_btb_made_pred;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_129 = T_38110_1_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_129 = T_38110_2_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_129 = T_38110_3_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_129 = T_38110_4_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_129 = T_38110_5_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_129 = T_38110_6_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_129 = T_38110_7_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_129 = T_38110_8_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_129 = T_38110_9_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_129 = T_38110_10_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_129 = T_38110_11_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_129 = T_38110_12_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_129 = T_38110_13_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_129 = T_38110_14_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_129 = T_38110_15_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_129 = T_38110_16_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_129 = T_38110_17_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_129 = T_38110_18_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_129 = T_38110_19_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_129 = T_38110_20_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_129 = T_38110_21_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_129 = T_38110_22_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_129 = T_38110_23_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_129 = T_38110_0_stat_btb_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_130 = T_38110_1_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_130 = T_38110_2_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_130 = T_38110_3_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_130 = T_38110_4_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_130 = T_38110_5_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_130 = T_38110_6_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_130 = T_38110_7_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_130 = T_38110_8_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_130 = T_38110_9_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_130 = T_38110_10_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_130 = T_38110_11_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_130 = T_38110_12_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_130 = T_38110_13_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_130 = T_38110_14_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_130 = T_38110_15_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_130 = T_38110_16_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_130 = T_38110_17_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_130 = T_38110_18_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_130 = T_38110_19_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_130 = T_38110_20_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_130 = T_38110_21_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_130 = T_38110_22_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_130 = T_38110_23_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_130 = T_38110_0_stat_bpd_made_pred;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_131 = T_38110_1_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_131 = T_38110_2_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_131 = T_38110_3_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_131 = T_38110_4_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_131 = T_38110_5_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_131 = T_38110_6_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_131 = T_38110_7_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_131 = T_38110_8_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_131 = T_38110_9_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_131 = T_38110_10_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_131 = T_38110_11_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_131 = T_38110_12_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_131 = T_38110_13_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_131 = T_38110_14_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_131 = T_38110_15_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_131 = T_38110_16_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_131 = T_38110_17_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_131 = T_38110_18_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_131 = T_38110_19_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_131 = T_38110_20_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_131 = T_38110_21_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_131 = T_38110_22_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_131 = T_38110_23_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_131 = T_38110_0_stat_bpd_mispredicted;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_132 = T_38110_1_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_132 = T_38110_2_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_132 = T_38110_3_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_132 = T_38110_4_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_132 = T_38110_5_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_132 = T_38110_6_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_132 = T_38110_7_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_132 = T_38110_8_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_132 = T_38110_9_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_132 = T_38110_10_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_132 = T_38110_11_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_132 = T_38110_12_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_132 = T_38110_13_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_132 = T_38110_14_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_132 = T_38110_15_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_132 = T_38110_16_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_132 = T_38110_17_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_132 = T_38110_18_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_132 = T_38110_19_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_132 = T_38110_20_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_132 = T_38110_21_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_132 = T_38110_22_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_132 = T_38110_23_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_132 = T_38110_0_fetch_pc_lob;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_133 = T_38110_1_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_133 = T_38110_2_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_133 = T_38110_3_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_133 = T_38110_4_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_133 = T_38110_5_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_133 = T_38110_6_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_133 = T_38110_7_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_133 = T_38110_8_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_133 = T_38110_9_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_133 = T_38110_10_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_133 = T_38110_11_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_133 = T_38110_12_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_133 = T_38110_13_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_133 = T_38110_14_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_133 = T_38110_15_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_133 = T_38110_16_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_133 = T_38110_17_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_133 = T_38110_18_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_133 = T_38110_19_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_133 = T_38110_20_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_133 = T_38110_21_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_133 = T_38110_22_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_133 = T_38110_23_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_133 = T_38110_0_imm_packed;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_134 = T_38110_1_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_134 = T_38110_2_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_134 = T_38110_3_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_134 = T_38110_4_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_134 = T_38110_5_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_134 = T_38110_6_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_134 = T_38110_7_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_134 = T_38110_8_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_134 = T_38110_9_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_134 = T_38110_10_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_134 = T_38110_11_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_134 = T_38110_12_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_134 = T_38110_13_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_134 = T_38110_14_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_134 = T_38110_15_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_134 = T_38110_16_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_134 = T_38110_17_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_134 = T_38110_18_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_134 = T_38110_19_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_134 = T_38110_20_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_134 = T_38110_21_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_134 = T_38110_22_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_134 = T_38110_23_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_134 = T_38110_0_csr_addr;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_135 = T_38110_1_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_135 = T_38110_2_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_135 = T_38110_3_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_135 = T_38110_4_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_135 = T_38110_5_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_135 = T_38110_6_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_135 = T_38110_7_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_135 = T_38110_8_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_135 = T_38110_9_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_135 = T_38110_10_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_135 = T_38110_11_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_135 = T_38110_12_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_135 = T_38110_13_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_135 = T_38110_14_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_135 = T_38110_15_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_135 = T_38110_16_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_135 = T_38110_17_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_135 = T_38110_18_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_135 = T_38110_19_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_135 = T_38110_20_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_135 = T_38110_21_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_135 = T_38110_22_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_135 = T_38110_23_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_135 = T_38110_0_rob_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_136 = T_38110_1_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_136 = T_38110_2_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_136 = T_38110_3_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_136 = T_38110_4_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_136 = T_38110_5_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_136 = T_38110_6_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_136 = T_38110_7_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_136 = T_38110_8_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_136 = T_38110_9_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_136 = T_38110_10_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_136 = T_38110_11_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_136 = T_38110_12_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_136 = T_38110_13_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_136 = T_38110_14_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_136 = T_38110_15_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_136 = T_38110_16_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_136 = T_38110_17_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_136 = T_38110_18_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_136 = T_38110_19_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_136 = T_38110_20_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_136 = T_38110_21_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_136 = T_38110_22_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_136 = T_38110_23_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_136 = T_38110_0_ldq_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_137 = T_38110_1_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_137 = T_38110_2_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_137 = T_38110_3_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_137 = T_38110_4_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_137 = T_38110_5_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_137 = T_38110_6_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_137 = T_38110_7_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_137 = T_38110_8_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_137 = T_38110_9_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_137 = T_38110_10_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_137 = T_38110_11_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_137 = T_38110_12_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_137 = T_38110_13_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_137 = T_38110_14_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_137 = T_38110_15_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_137 = T_38110_16_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_137 = T_38110_17_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_137 = T_38110_18_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_137 = T_38110_19_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_137 = T_38110_20_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_137 = T_38110_21_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_137 = T_38110_22_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_137 = T_38110_23_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_137 = T_38110_0_stq_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_138 = T_38110_1_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_138 = T_38110_2_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_138 = T_38110_3_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_138 = T_38110_4_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_138 = T_38110_5_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_138 = T_38110_6_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_138 = T_38110_7_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_138 = T_38110_8_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_138 = T_38110_9_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_138 = T_38110_10_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_138 = T_38110_11_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_138 = T_38110_12_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_138 = T_38110_13_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_138 = T_38110_14_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_138 = T_38110_15_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_138 = T_38110_16_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_138 = T_38110_17_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_138 = T_38110_18_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_138 = T_38110_19_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_138 = T_38110_20_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_138 = T_38110_21_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_138 = T_38110_22_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_138 = T_38110_23_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_138 = T_38110_0_brob_idx;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_139 = T_38110_1_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_139 = T_38110_2_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_139 = T_38110_3_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_139 = T_38110_4_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_139 = T_38110_5_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_139 = T_38110_6_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_139 = T_38110_7_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_139 = T_38110_8_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_139 = T_38110_9_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_139 = T_38110_10_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_139 = T_38110_11_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_139 = T_38110_12_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_139 = T_38110_13_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_139 = T_38110_14_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_139 = T_38110_15_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_139 = T_38110_16_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_139 = T_38110_17_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_139 = T_38110_18_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_139 = T_38110_19_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_139 = T_38110_20_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_139 = T_38110_21_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_139 = T_38110_22_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_139 = T_38110_23_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_139 = T_38110_0_pdst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_140 = T_38110_1_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_140 = T_38110_2_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_140 = T_38110_3_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_140 = T_38110_4_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_140 = T_38110_5_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_140 = T_38110_6_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_140 = T_38110_7_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_140 = T_38110_8_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_140 = T_38110_9_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_140 = T_38110_10_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_140 = T_38110_11_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_140 = T_38110_12_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_140 = T_38110_13_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_140 = T_38110_14_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_140 = T_38110_15_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_140 = T_38110_16_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_140 = T_38110_17_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_140 = T_38110_18_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_140 = T_38110_19_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_140 = T_38110_20_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_140 = T_38110_21_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_140 = T_38110_22_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_140 = T_38110_23_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_140 = T_38110_0_pop1;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_141 = T_38110_1_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_141 = T_38110_2_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_141 = T_38110_3_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_141 = T_38110_4_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_141 = T_38110_5_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_141 = T_38110_6_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_141 = T_38110_7_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_141 = T_38110_8_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_141 = T_38110_9_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_141 = T_38110_10_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_141 = T_38110_11_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_141 = T_38110_12_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_141 = T_38110_13_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_141 = T_38110_14_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_141 = T_38110_15_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_141 = T_38110_16_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_141 = T_38110_17_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_141 = T_38110_18_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_141 = T_38110_19_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_141 = T_38110_20_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_141 = T_38110_21_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_141 = T_38110_22_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_141 = T_38110_23_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_141 = T_38110_0_pop2;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_142 = T_38110_1_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_142 = T_38110_2_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_142 = T_38110_3_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_142 = T_38110_4_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_142 = T_38110_5_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_142 = T_38110_6_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_142 = T_38110_7_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_142 = T_38110_8_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_142 = T_38110_9_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_142 = T_38110_10_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_142 = T_38110_11_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_142 = T_38110_12_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_142 = T_38110_13_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_142 = T_38110_14_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_142 = T_38110_15_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_142 = T_38110_16_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_142 = T_38110_17_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_142 = T_38110_18_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_142 = T_38110_19_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_142 = T_38110_20_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_142 = T_38110_21_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_142 = T_38110_22_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_142 = T_38110_23_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_142 = T_38110_0_pop3;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_143 = T_38110_1_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_143 = T_38110_2_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_143 = T_38110_3_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_143 = T_38110_4_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_143 = T_38110_5_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_143 = T_38110_6_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_143 = T_38110_7_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_143 = T_38110_8_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_143 = T_38110_9_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_143 = T_38110_10_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_143 = T_38110_11_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_143 = T_38110_12_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_143 = T_38110_13_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_143 = T_38110_14_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_143 = T_38110_15_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_143 = T_38110_16_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_143 = T_38110_17_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_143 = T_38110_18_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_143 = T_38110_19_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_143 = T_38110_20_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_143 = T_38110_21_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_143 = T_38110_22_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_143 = T_38110_23_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_143 = T_38110_0_prs1_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_144 = T_38110_1_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_144 = T_38110_2_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_144 = T_38110_3_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_144 = T_38110_4_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_144 = T_38110_5_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_144 = T_38110_6_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_144 = T_38110_7_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_144 = T_38110_8_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_144 = T_38110_9_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_144 = T_38110_10_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_144 = T_38110_11_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_144 = T_38110_12_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_144 = T_38110_13_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_144 = T_38110_14_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_144 = T_38110_15_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_144 = T_38110_16_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_144 = T_38110_17_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_144 = T_38110_18_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_144 = T_38110_19_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_144 = T_38110_20_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_144 = T_38110_21_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_144 = T_38110_22_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_144 = T_38110_23_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_144 = T_38110_0_prs2_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_145 = T_38110_1_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_145 = T_38110_2_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_145 = T_38110_3_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_145 = T_38110_4_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_145 = T_38110_5_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_145 = T_38110_6_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_145 = T_38110_7_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_145 = T_38110_8_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_145 = T_38110_9_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_145 = T_38110_10_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_145 = T_38110_11_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_145 = T_38110_12_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_145 = T_38110_13_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_145 = T_38110_14_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_145 = T_38110_15_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_145 = T_38110_16_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_145 = T_38110_17_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_145 = T_38110_18_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_145 = T_38110_19_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_145 = T_38110_20_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_145 = T_38110_21_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_145 = T_38110_22_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_145 = T_38110_23_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_145 = T_38110_0_prs3_busy;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_146 = T_38110_1_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_146 = T_38110_2_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_146 = T_38110_3_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_146 = T_38110_4_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_146 = T_38110_5_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_146 = T_38110_6_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_146 = T_38110_7_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_146 = T_38110_8_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_146 = T_38110_9_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_146 = T_38110_10_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_146 = T_38110_11_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_146 = T_38110_12_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_146 = T_38110_13_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_146 = T_38110_14_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_146 = T_38110_15_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_146 = T_38110_16_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_146 = T_38110_17_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_146 = T_38110_18_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_146 = T_38110_19_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_146 = T_38110_20_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_146 = T_38110_21_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_146 = T_38110_22_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_146 = T_38110_23_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_146 = T_38110_0_stale_pdst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_147 = T_38110_1_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_147 = T_38110_2_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_147 = T_38110_3_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_147 = T_38110_4_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_147 = T_38110_5_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_147 = T_38110_6_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_147 = T_38110_7_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_147 = T_38110_8_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_147 = T_38110_9_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_147 = T_38110_10_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_147 = T_38110_11_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_147 = T_38110_12_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_147 = T_38110_13_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_147 = T_38110_14_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_147 = T_38110_15_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_147 = T_38110_16_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_147 = T_38110_17_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_147 = T_38110_18_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_147 = T_38110_19_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_147 = T_38110_20_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_147 = T_38110_21_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_147 = T_38110_22_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_147 = T_38110_23_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_147 = T_38110_0_exception;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_148 = T_38110_1_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_148 = T_38110_2_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_148 = T_38110_3_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_148 = T_38110_4_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_148 = T_38110_5_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_148 = T_38110_6_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_148 = T_38110_7_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_148 = T_38110_8_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_148 = T_38110_9_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_148 = T_38110_10_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_148 = T_38110_11_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_148 = T_38110_12_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_148 = T_38110_13_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_148 = T_38110_14_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_148 = T_38110_15_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_148 = T_38110_16_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_148 = T_38110_17_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_148 = T_38110_18_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_148 = T_38110_19_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_148 = T_38110_20_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_148 = T_38110_21_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_148 = T_38110_22_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_148 = T_38110_23_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_148 = T_38110_0_exc_cause;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_149 = T_38110_1_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_149 = T_38110_2_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_149 = T_38110_3_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_149 = T_38110_4_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_149 = T_38110_5_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_149 = T_38110_6_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_149 = T_38110_7_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_149 = T_38110_8_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_149 = T_38110_9_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_149 = T_38110_10_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_149 = T_38110_11_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_149 = T_38110_12_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_149 = T_38110_13_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_149 = T_38110_14_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_149 = T_38110_15_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_149 = T_38110_16_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_149 = T_38110_17_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_149 = T_38110_18_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_149 = T_38110_19_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_149 = T_38110_20_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_149 = T_38110_21_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_149 = T_38110_22_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_149 = T_38110_23_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_149 = T_38110_0_bypassable;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_150 = T_38110_1_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_150 = T_38110_2_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_150 = T_38110_3_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_150 = T_38110_4_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_150 = T_38110_5_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_150 = T_38110_6_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_150 = T_38110_7_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_150 = T_38110_8_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_150 = T_38110_9_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_150 = T_38110_10_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_150 = T_38110_11_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_150 = T_38110_12_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_150 = T_38110_13_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_150 = T_38110_14_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_150 = T_38110_15_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_150 = T_38110_16_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_150 = T_38110_17_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_150 = T_38110_18_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_150 = T_38110_19_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_150 = T_38110_20_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_150 = T_38110_21_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_150 = T_38110_22_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_150 = T_38110_23_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_150 = T_38110_0_mem_cmd;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_151 = T_38110_1_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_151 = T_38110_2_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_151 = T_38110_3_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_151 = T_38110_4_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_151 = T_38110_5_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_151 = T_38110_6_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_151 = T_38110_7_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_151 = T_38110_8_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_151 = T_38110_9_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_151 = T_38110_10_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_151 = T_38110_11_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_151 = T_38110_12_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_151 = T_38110_13_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_151 = T_38110_14_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_151 = T_38110_15_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_151 = T_38110_16_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_151 = T_38110_17_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_151 = T_38110_18_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_151 = T_38110_19_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_151 = T_38110_20_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_151 = T_38110_21_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_151 = T_38110_22_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_151 = T_38110_23_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_151 = T_38110_0_mem_typ;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_152 = T_38110_1_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_152 = T_38110_2_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_152 = T_38110_3_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_152 = T_38110_4_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_152 = T_38110_5_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_152 = T_38110_6_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_152 = T_38110_7_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_152 = T_38110_8_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_152 = T_38110_9_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_152 = T_38110_10_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_152 = T_38110_11_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_152 = T_38110_12_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_152 = T_38110_13_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_152 = T_38110_14_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_152 = T_38110_15_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_152 = T_38110_16_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_152 = T_38110_17_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_152 = T_38110_18_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_152 = T_38110_19_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_152 = T_38110_20_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_152 = T_38110_21_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_152 = T_38110_22_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_152 = T_38110_23_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_152 = T_38110_0_is_fence;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_153 = T_38110_1_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_153 = T_38110_2_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_153 = T_38110_3_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_153 = T_38110_4_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_153 = T_38110_5_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_153 = T_38110_6_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_153 = T_38110_7_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_153 = T_38110_8_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_153 = T_38110_9_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_153 = T_38110_10_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_153 = T_38110_11_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_153 = T_38110_12_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_153 = T_38110_13_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_153 = T_38110_14_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_153 = T_38110_15_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_153 = T_38110_16_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_153 = T_38110_17_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_153 = T_38110_18_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_153 = T_38110_19_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_153 = T_38110_20_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_153 = T_38110_21_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_153 = T_38110_22_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_153 = T_38110_23_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_153 = T_38110_0_is_fencei;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_154 = T_38110_1_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_154 = T_38110_2_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_154 = T_38110_3_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_154 = T_38110_4_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_154 = T_38110_5_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_154 = T_38110_6_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_154 = T_38110_7_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_154 = T_38110_8_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_154 = T_38110_9_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_154 = T_38110_10_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_154 = T_38110_11_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_154 = T_38110_12_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_154 = T_38110_13_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_154 = T_38110_14_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_154 = T_38110_15_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_154 = T_38110_16_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_154 = T_38110_17_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_154 = T_38110_18_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_154 = T_38110_19_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_154 = T_38110_20_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_154 = T_38110_21_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_154 = T_38110_22_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_154 = T_38110_23_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_154 = T_38110_0_is_store;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_155 = T_38110_1_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_155 = T_38110_2_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_155 = T_38110_3_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_155 = T_38110_4_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_155 = T_38110_5_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_155 = T_38110_6_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_155 = T_38110_7_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_155 = T_38110_8_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_155 = T_38110_9_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_155 = T_38110_10_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_155 = T_38110_11_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_155 = T_38110_12_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_155 = T_38110_13_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_155 = T_38110_14_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_155 = T_38110_15_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_155 = T_38110_16_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_155 = T_38110_17_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_155 = T_38110_18_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_155 = T_38110_19_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_155 = T_38110_20_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_155 = T_38110_21_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_155 = T_38110_22_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_155 = T_38110_23_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_155 = T_38110_0_is_amo;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_156 = T_38110_1_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_156 = T_38110_2_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_156 = T_38110_3_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_156 = T_38110_4_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_156 = T_38110_5_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_156 = T_38110_6_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_156 = T_38110_7_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_156 = T_38110_8_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_156 = T_38110_9_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_156 = T_38110_10_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_156 = T_38110_11_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_156 = T_38110_12_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_156 = T_38110_13_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_156 = T_38110_14_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_156 = T_38110_15_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_156 = T_38110_16_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_156 = T_38110_17_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_156 = T_38110_18_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_156 = T_38110_19_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_156 = T_38110_20_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_156 = T_38110_21_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_156 = T_38110_22_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_156 = T_38110_23_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_156 = T_38110_0_is_load;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_157 = T_38110_1_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_157 = T_38110_2_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_157 = T_38110_3_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_157 = T_38110_4_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_157 = T_38110_5_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_157 = T_38110_6_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_157 = T_38110_7_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_157 = T_38110_8_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_157 = T_38110_9_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_157 = T_38110_10_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_157 = T_38110_11_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_157 = T_38110_12_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_157 = T_38110_13_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_157 = T_38110_14_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_157 = T_38110_15_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_157 = T_38110_16_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_157 = T_38110_17_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_157 = T_38110_18_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_157 = T_38110_19_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_157 = T_38110_20_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_157 = T_38110_21_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_157 = T_38110_22_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_157 = T_38110_23_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_157 = T_38110_0_is_unique;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_158 = T_38110_1_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_158 = T_38110_2_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_158 = T_38110_3_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_158 = T_38110_4_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_158 = T_38110_5_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_158 = T_38110_6_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_158 = T_38110_7_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_158 = T_38110_8_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_158 = T_38110_9_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_158 = T_38110_10_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_158 = T_38110_11_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_158 = T_38110_12_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_158 = T_38110_13_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_158 = T_38110_14_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_158 = T_38110_15_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_158 = T_38110_16_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_158 = T_38110_17_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_158 = T_38110_18_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_158 = T_38110_19_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_158 = T_38110_20_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_158 = T_38110_21_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_158 = T_38110_22_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_158 = T_38110_23_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_158 = T_38110_0_flush_on_commit;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_159 = T_38110_1_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_159 = T_38110_2_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_159 = T_38110_3_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_159 = T_38110_4_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_159 = T_38110_5_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_159 = T_38110_6_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_159 = T_38110_7_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_159 = T_38110_8_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_159 = T_38110_9_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_159 = T_38110_10_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_159 = T_38110_11_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_159 = T_38110_12_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_159 = T_38110_13_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_159 = T_38110_14_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_159 = T_38110_15_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_159 = T_38110_16_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_159 = T_38110_17_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_159 = T_38110_18_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_159 = T_38110_19_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_159 = T_38110_20_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_159 = T_38110_21_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_159 = T_38110_22_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_159 = T_38110_23_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_159 = T_38110_0_ldst;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_160 = T_38110_1_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_160 = T_38110_2_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_160 = T_38110_3_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_160 = T_38110_4_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_160 = T_38110_5_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_160 = T_38110_6_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_160 = T_38110_7_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_160 = T_38110_8_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_160 = T_38110_9_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_160 = T_38110_10_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_160 = T_38110_11_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_160 = T_38110_12_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_160 = T_38110_13_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_160 = T_38110_14_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_160 = T_38110_15_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_160 = T_38110_16_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_160 = T_38110_17_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_160 = T_38110_18_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_160 = T_38110_19_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_160 = T_38110_20_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_160 = T_38110_21_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_160 = T_38110_22_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_160 = T_38110_23_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_160 = T_38110_0_lrs1;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_161 = T_38110_1_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_161 = T_38110_2_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_161 = T_38110_3_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_161 = T_38110_4_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_161 = T_38110_5_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_161 = T_38110_6_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_161 = T_38110_7_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_161 = T_38110_8_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_161 = T_38110_9_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_161 = T_38110_10_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_161 = T_38110_11_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_161 = T_38110_12_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_161 = T_38110_13_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_161 = T_38110_14_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_161 = T_38110_15_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_161 = T_38110_16_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_161 = T_38110_17_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_161 = T_38110_18_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_161 = T_38110_19_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_161 = T_38110_20_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_161 = T_38110_21_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_161 = T_38110_22_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_161 = T_38110_23_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_161 = T_38110_0_lrs2;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_162 = T_38110_1_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_162 = T_38110_2_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_162 = T_38110_3_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_162 = T_38110_4_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_162 = T_38110_5_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_162 = T_38110_6_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_162 = T_38110_7_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_162 = T_38110_8_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_162 = T_38110_9_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_162 = T_38110_10_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_162 = T_38110_11_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_162 = T_38110_12_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_162 = T_38110_13_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_162 = T_38110_14_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_162 = T_38110_15_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_162 = T_38110_16_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_162 = T_38110_17_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_162 = T_38110_18_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_162 = T_38110_19_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_162 = T_38110_20_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_162 = T_38110_21_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_162 = T_38110_22_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_162 = T_38110_23_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_162 = T_38110_0_lrs3;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_163 = T_38110_1_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_163 = T_38110_2_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_163 = T_38110_3_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_163 = T_38110_4_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_163 = T_38110_5_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_163 = T_38110_6_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_163 = T_38110_7_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_163 = T_38110_8_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_163 = T_38110_9_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_163 = T_38110_10_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_163 = T_38110_11_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_163 = T_38110_12_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_163 = T_38110_13_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_163 = T_38110_14_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_163 = T_38110_15_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_163 = T_38110_16_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_163 = T_38110_17_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_163 = T_38110_18_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_163 = T_38110_19_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_163 = T_38110_20_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_163 = T_38110_21_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_163 = T_38110_22_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_163 = T_38110_23_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_163 = T_38110_0_ldst_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_164 = T_38110_1_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_164 = T_38110_2_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_164 = T_38110_3_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_164 = T_38110_4_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_164 = T_38110_5_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_164 = T_38110_6_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_164 = T_38110_7_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_164 = T_38110_8_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_164 = T_38110_9_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_164 = T_38110_10_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_164 = T_38110_11_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_164 = T_38110_12_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_164 = T_38110_13_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_164 = T_38110_14_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_164 = T_38110_15_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_164 = T_38110_16_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_164 = T_38110_17_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_164 = T_38110_18_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_164 = T_38110_19_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_164 = T_38110_20_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_164 = T_38110_21_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_164 = T_38110_22_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_164 = T_38110_23_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_164 = T_38110_0_dst_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_165 = T_38110_1_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_165 = T_38110_2_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_165 = T_38110_3_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_165 = T_38110_4_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_165 = T_38110_5_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_165 = T_38110_6_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_165 = T_38110_7_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_165 = T_38110_8_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_165 = T_38110_9_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_165 = T_38110_10_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_165 = T_38110_11_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_165 = T_38110_12_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_165 = T_38110_13_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_165 = T_38110_14_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_165 = T_38110_15_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_165 = T_38110_16_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_165 = T_38110_17_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_165 = T_38110_18_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_165 = T_38110_19_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_165 = T_38110_20_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_165 = T_38110_21_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_165 = T_38110_22_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_165 = T_38110_23_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_165 = T_38110_0_lrs1_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_166 = T_38110_1_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_166 = T_38110_2_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_166 = T_38110_3_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_166 = T_38110_4_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_166 = T_38110_5_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_166 = T_38110_6_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_166 = T_38110_7_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_166 = T_38110_8_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_166 = T_38110_9_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_166 = T_38110_10_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_166 = T_38110_11_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_166 = T_38110_12_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_166 = T_38110_13_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_166 = T_38110_14_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_166 = T_38110_15_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_166 = T_38110_16_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_166 = T_38110_17_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_166 = T_38110_18_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_166 = T_38110_19_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_166 = T_38110_20_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_166 = T_38110_21_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_166 = T_38110_22_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_166 = T_38110_23_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_166 = T_38110_0_lrs2_rtype;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_167 = T_38110_1_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_167 = T_38110_2_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_167 = T_38110_3_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_167 = T_38110_4_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_167 = T_38110_5_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_167 = T_38110_6_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_167 = T_38110_7_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_167 = T_38110_8_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_167 = T_38110_9_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_167 = T_38110_10_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_167 = T_38110_11_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_167 = T_38110_12_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_167 = T_38110_13_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_167 = T_38110_14_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_167 = T_38110_15_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_167 = T_38110_16_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_167 = T_38110_17_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_167 = T_38110_18_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_167 = T_38110_19_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_167 = T_38110_20_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_167 = T_38110_21_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_167 = T_38110_22_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_167 = T_38110_23_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_167 = T_38110_0_frs3_en;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_168 = T_38110_1_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_168 = T_38110_2_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_168 = T_38110_3_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_168 = T_38110_4_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_168 = T_38110_5_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_168 = T_38110_6_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_168 = T_38110_7_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_168 = T_38110_8_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_168 = T_38110_9_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_168 = T_38110_10_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_168 = T_38110_11_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_168 = T_38110_12_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_168 = T_38110_13_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_168 = T_38110_14_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_168 = T_38110_15_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_168 = T_38110_16_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_168 = T_38110_17_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_168 = T_38110_18_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_168 = T_38110_19_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_168 = T_38110_20_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_168 = T_38110_21_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_168 = T_38110_22_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_168 = T_38110_23_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_168 = T_38110_0_fp_val;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_169 = T_38110_1_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_169 = T_38110_2_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_169 = T_38110_3_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_169 = T_38110_4_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_169 = T_38110_5_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_169 = T_38110_6_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_169 = T_38110_7_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_169 = T_38110_8_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_169 = T_38110_9_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_169 = T_38110_10_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_169 = T_38110_11_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_169 = T_38110_12_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_169 = T_38110_13_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_169 = T_38110_14_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_169 = T_38110_15_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_169 = T_38110_16_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_169 = T_38110_17_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_169 = T_38110_18_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_169 = T_38110_19_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_169 = T_38110_20_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_169 = T_38110_21_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_169 = T_38110_22_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_169 = T_38110_23_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_169 = T_38110_0_fp_single;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_170 = T_38110_1_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_170 = T_38110_2_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_170 = T_38110_3_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_170 = T_38110_4_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_170 = T_38110_5_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_170 = T_38110_6_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_170 = T_38110_7_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_170 = T_38110_8_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_170 = T_38110_9_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_170 = T_38110_10_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_170 = T_38110_11_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_170 = T_38110_12_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_170 = T_38110_13_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_170 = T_38110_14_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_170 = T_38110_15_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_170 = T_38110_16_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_170 = T_38110_17_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_170 = T_38110_18_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_170 = T_38110_19_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_170 = T_38110_20_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_170 = T_38110_21_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_170 = T_38110_22_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_170 = T_38110_23_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_170 = T_38110_0_xcpt_if;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_171 = T_38110_1_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_171 = T_38110_2_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_171 = T_38110_3_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_171 = T_38110_4_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_171 = T_38110_5_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_171 = T_38110_6_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_171 = T_38110_7_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_171 = T_38110_8_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_171 = T_38110_9_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_171 = T_38110_10_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_171 = T_38110_11_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_171 = T_38110_12_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_171 = T_38110_13_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_171 = T_38110_14_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_171 = T_38110_15_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_171 = T_38110_16_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_171 = T_38110_17_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_171 = T_38110_18_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_171 = T_38110_19_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_171 = T_38110_20_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_171 = T_38110_21_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_171 = T_38110_22_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_171 = T_38110_23_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_171 = T_38110_0_replay_if;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:451:58, :453:59
    casez (_T_2)	// rob.scala:451:58, :453:59
      5'b00000:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00001:
        casez_tmp_172 = T_38110_1_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00010:
        casez_tmp_172 = T_38110_2_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00011:
        casez_tmp_172 = T_38110_3_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00100:
        casez_tmp_172 = T_38110_4_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00101:
        casez_tmp_172 = T_38110_5_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00110:
        casez_tmp_172 = T_38110_6_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b00111:
        casez_tmp_172 = T_38110_7_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01000:
        casez_tmp_172 = T_38110_8_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01001:
        casez_tmp_172 = T_38110_9_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01010:
        casez_tmp_172 = T_38110_10_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01011:
        casez_tmp_172 = T_38110_11_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01100:
        casez_tmp_172 = T_38110_12_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01101:
        casez_tmp_172 = T_38110_13_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01110:
        casez_tmp_172 = T_38110_14_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b01111:
        casez_tmp_172 = T_38110_15_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10000:
        casez_tmp_172 = T_38110_16_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10001:
        casez_tmp_172 = T_38110_17_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10010:
        casez_tmp_172 = T_38110_18_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10011:
        casez_tmp_172 = T_38110_19_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10100:
        casez_tmp_172 = T_38110_20_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10101:
        casez_tmp_172 = T_38110_21_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10110:
        casez_tmp_172 = T_38110_22_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b10111:
        casez_tmp_172 = T_38110_23_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11000:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11001:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11010:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11011:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11100:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11101:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      5'b11110:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
      default:
        casez_tmp_172 = T_38110_0_debug_events_fetch_seq;	// rob.scala:350:34, :451:58, :453:59
    endcase	// rob.scala:451:58, :453:59
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_173 = T_38110_1_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_173 = T_38110_2_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_173 = T_38110_3_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_173 = T_38110_4_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_173 = T_38110_5_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_173 = T_38110_6_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_173 = T_38110_7_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_173 = T_38110_8_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_173 = T_38110_9_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_173 = T_38110_10_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_173 = T_38110_11_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_173 = T_38110_12_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_173 = T_38110_13_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_173 = T_38110_14_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_173 = T_38110_15_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_173 = T_38110_16_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_173 = T_38110_17_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_173 = T_38110_18_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_173 = T_38110_19_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_173 = T_38110_20_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_173 = T_38110_21_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_173 = T_38110_22_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_173 = T_38110_23_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_173 = T_38110_0_is_store;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_174 = T_38110_1_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_174 = T_38110_2_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_174 = T_38110_3_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_174 = T_38110_4_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_174 = T_38110_5_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_174 = T_38110_6_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_174 = T_38110_7_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_174 = T_38110_8_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_174 = T_38110_9_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_174 = T_38110_10_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_174 = T_38110_11_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_174 = T_38110_12_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_174 = T_38110_13_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_174 = T_38110_14_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_174 = T_38110_15_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_174 = T_38110_16_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_174 = T_38110_17_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_174 = T_38110_18_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_174 = T_38110_19_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_174 = T_38110_20_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_174 = T_38110_21_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_174 = T_38110_22_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_174 = T_38110_23_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_174 = T_38110_0_is_load;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  always @(*) begin	// rob.scala:433:51, :507:28
    casez (rob_head)	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
      5'b00000:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00001:
        casez_tmp_175 = T_38110_1_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00010:
        casez_tmp_175 = T_38110_2_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00011:
        casez_tmp_175 = T_38110_3_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00100:
        casez_tmp_175 = T_38110_4_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00101:
        casez_tmp_175 = T_38110_5_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00110:
        casez_tmp_175 = T_38110_6_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b00111:
        casez_tmp_175 = T_38110_7_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01000:
        casez_tmp_175 = T_38110_8_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01001:
        casez_tmp_175 = T_38110_9_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01010:
        casez_tmp_175 = T_38110_10_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01011:
        casez_tmp_175 = T_38110_11_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01100:
        casez_tmp_175 = T_38110_12_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01101:
        casez_tmp_175 = T_38110_13_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01110:
        casez_tmp_175 = T_38110_14_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b01111:
        casez_tmp_175 = T_38110_15_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10000:
        casez_tmp_175 = T_38110_16_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10001:
        casez_tmp_175 = T_38110_17_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10010:
        casez_tmp_175 = T_38110_18_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10011:
        casez_tmp_175 = T_38110_19_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10100:
        casez_tmp_175 = T_38110_20_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10101:
        casez_tmp_175 = T_38110_21_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10110:
        casez_tmp_175 = T_38110_22_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b10111:
        casez_tmp_175 = T_38110_23_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11000:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11001:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11010:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11011:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11100:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11101:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      5'b11110:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
      default:
        casez_tmp_175 = T_38110_0_debug_wdata;	// rob.scala:350:34, :433:51, :507:28
    endcase	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:433:51, :507:28
  end // always @(*)
  wire [5:0] _T_43921 = _io_get_pc_rob_idx_5to1 == 5'h17 ? 6'h0 : {1'h0, _io_get_pc_rob_idx_5to1} + 6'h1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:347:34, :967:16, util.scala:75:28, :76:{13,35}
  assign _T_0 = _T_43921 == 6'h17 ? T_35634_23 : _T_43921 == 6'h16 ? T_35634_22 : _T_43921 == 6'h15 ?
                T_35634_21 : _T_43921 == 6'h14 ? T_35634_20 : _T_43921 == 6'h13 ? T_35634_19 : _T_43921 ==
                6'h12 ? T_35634_18 : _T_43921 == 6'h11 ? T_35634_17 : _T_43921 == 6'h10 ? T_35634_16 :
                _T_43921 == 6'hF ? T_35634_15 : _T_43921 == 6'hE ? T_35634_14 : _T_43921 == 6'hD ?
                T_35634_13 : _T_43921 == 6'hC ? T_35634_12 : _T_43921 == 6'hB ? T_35634_11 : _T_43921 ==
                6'hA ? T_35634_10 : _T_43921 == 6'h9 ? T_35634_9 : _T_43921 == 6'h8 ? T_35634_8 : _T_43921
                == 6'h7 ? T_35634_7 : _T_43921 == 6'h6 ? T_35634_6 : _T_43921 == 6'h5 ? T_35634_5 :
                _T_43921 == 6'h4 ? T_35634_4 : _T_43921 == 6'h3 ? T_35634_3 : _T_43921 == 6'h2 ? T_35634_2
                : _T_43921 == 6'h1 ? T_35634_1 : T_35634_0;	// rob.scala:347:34, :509:28, :967:16
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_176 = T_35634_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_176 = T_35634_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_176 = T_35634_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_176 = T_35634_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_176 = T_35634_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_176 = T_35634_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_176 = T_35634_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_176 = T_35634_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_176 = T_35634_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_176 = T_35634_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_176 = T_35634_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_176 = T_35634_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_176 = T_35634_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_176 = T_35634_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_176 = T_35634_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_176 = T_35634_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_176 = T_35634_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_176 = T_35634_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_176 = T_35634_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_176 = T_35634_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_176 = T_35634_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_176 = T_35634_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_176 = T_35634_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_176 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_177 = T_38110_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_177 = T_38110_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_177 = T_38110_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_177 = T_38110_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_177 = T_38110_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_177 = T_38110_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_177 = T_38110_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_177 = T_38110_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_177 = T_38110_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_177 = T_38110_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_177 = T_38110_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_177 = T_38110_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_177 = T_38110_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_177 = T_38110_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_177 = T_38110_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_177 = T_38110_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_177 = T_38110_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_177 = T_38110_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_177 = T_38110_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_177 = T_38110_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_177 = T_38110_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_177 = T_38110_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_177 = T_38110_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_177 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_0_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_178 = T_38110_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_178 = T_38110_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_178 = T_38110_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_178 = T_38110_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_178 = T_38110_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_178 = T_38110_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_178 = T_38110_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_178 = T_38110_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_178 = T_38110_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_178 = T_38110_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_178 = T_38110_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_178 = T_38110_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_178 = T_38110_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_178 = T_38110_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_178 = T_38110_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_178 = T_38110_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_178 = T_38110_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_178 = T_38110_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_178 = T_38110_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_178 = T_38110_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_178 = T_38110_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_178 = T_38110_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_178 = T_38110_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_178 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_179 = T_35634_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_179 = T_35634_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_179 = T_35634_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_179 = T_35634_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_179 = T_35634_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_179 = T_35634_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_179 = T_35634_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_179 = T_35634_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_179 = T_35634_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_179 = T_35634_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_179 = T_35634_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_179 = T_35634_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_179 = T_35634_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_179 = T_35634_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_179 = T_35634_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_179 = T_35634_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_179 = T_35634_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_179 = T_35634_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_179 = T_35634_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_179 = T_35634_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_179 = T_35634_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_179 = T_35634_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_179 = T_35634_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_179 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_180 = T_38110_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_180 = T_38110_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_180 = T_38110_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_180 = T_38110_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_180 = T_38110_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_180 = T_38110_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_180 = T_38110_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_180 = T_38110_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_180 = T_38110_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_180 = T_38110_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_180 = T_38110_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_180 = T_38110_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_180 = T_38110_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_180 = T_38110_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_180 = T_38110_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_180 = T_38110_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_180 = T_38110_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_180 = T_38110_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_180 = T_38110_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_180 = T_38110_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_180 = T_38110_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_180 = T_38110_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_180 = T_38110_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_180 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_1_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_181 = T_38110_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_181 = T_38110_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_181 = T_38110_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_181 = T_38110_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_181 = T_38110_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_181 = T_38110_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_181 = T_38110_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_181 = T_38110_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_181 = T_38110_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_181 = T_38110_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_181 = T_38110_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_181 = T_38110_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_181 = T_38110_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_181 = T_38110_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_181 = T_38110_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_181 = T_38110_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_181 = T_38110_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_181 = T_38110_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_181 = T_38110_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_181 = T_38110_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_181 = T_38110_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_181 = T_38110_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_181 = T_38110_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_181 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :536:22
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :536:22
      5'b00000:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b00001:
        casez_tmp_182 = T_35634_1;	// rob.scala:347:34, :531:53, :536:22
      5'b00010:
        casez_tmp_182 = T_35634_2;	// rob.scala:347:34, :531:53, :536:22
      5'b00011:
        casez_tmp_182 = T_35634_3;	// rob.scala:347:34, :531:53, :536:22
      5'b00100:
        casez_tmp_182 = T_35634_4;	// rob.scala:347:34, :531:53, :536:22
      5'b00101:
        casez_tmp_182 = T_35634_5;	// rob.scala:347:34, :531:53, :536:22
      5'b00110:
        casez_tmp_182 = T_35634_6;	// rob.scala:347:34, :531:53, :536:22
      5'b00111:
        casez_tmp_182 = T_35634_7;	// rob.scala:347:34, :531:53, :536:22
      5'b01000:
        casez_tmp_182 = T_35634_8;	// rob.scala:347:34, :531:53, :536:22
      5'b01001:
        casez_tmp_182 = T_35634_9;	// rob.scala:347:34, :531:53, :536:22
      5'b01010:
        casez_tmp_182 = T_35634_10;	// rob.scala:347:34, :531:53, :536:22
      5'b01011:
        casez_tmp_182 = T_35634_11;	// rob.scala:347:34, :531:53, :536:22
      5'b01100:
        casez_tmp_182 = T_35634_12;	// rob.scala:347:34, :531:53, :536:22
      5'b01101:
        casez_tmp_182 = T_35634_13;	// rob.scala:347:34, :531:53, :536:22
      5'b01110:
        casez_tmp_182 = T_35634_14;	// rob.scala:347:34, :531:53, :536:22
      5'b01111:
        casez_tmp_182 = T_35634_15;	// rob.scala:347:34, :531:53, :536:22
      5'b10000:
        casez_tmp_182 = T_35634_16;	// rob.scala:347:34, :531:53, :536:22
      5'b10001:
        casez_tmp_182 = T_35634_17;	// rob.scala:347:34, :531:53, :536:22
      5'b10010:
        casez_tmp_182 = T_35634_18;	// rob.scala:347:34, :531:53, :536:22
      5'b10011:
        casez_tmp_182 = T_35634_19;	// rob.scala:347:34, :531:53, :536:22
      5'b10100:
        casez_tmp_182 = T_35634_20;	// rob.scala:347:34, :531:53, :536:22
      5'b10101:
        casez_tmp_182 = T_35634_21;	// rob.scala:347:34, :531:53, :536:22
      5'b10110:
        casez_tmp_182 = T_35634_22;	// rob.scala:347:34, :531:53, :536:22
      5'b10111:
        casez_tmp_182 = T_35634_23;	// rob.scala:347:34, :531:53, :536:22
      5'b11000:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11001:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11010:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11011:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11100:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11101:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      5'b11110:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
      default:
        casez_tmp_182 = T_35634_0;	// rob.scala:347:34, :531:53, :536:22
    endcase	// rob.scala:531:53, :536:22
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_183 = T_38110_1_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_183 = T_38110_2_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_183 = T_38110_3_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_183 = T_38110_4_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_183 = T_38110_5_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_183 = T_38110_6_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_183 = T_38110_7_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_183 = T_38110_8_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_183 = T_38110_9_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_183 = T_38110_10_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_183 = T_38110_11_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_183 = T_38110_12_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_183 = T_38110_13_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_183 = T_38110_14_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_183 = T_38110_15_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_183 = T_38110_16_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_183 = T_38110_17_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_183 = T_38110_18_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_183 = T_38110_19_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_183 = T_38110_20_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_183 = T_38110_21_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_183 = T_38110_22_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_183 = T_38110_23_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_183 = T_38110_0_pdst;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  always @(*) begin	// rob.scala:531:53, :538:75
    casez (_io_wb_resps_2_bits_uop_rob_idx_5to1)	// rob.scala:531:53, :538:75
      5'b00000:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00001:
        casez_tmp_184 = T_38110_1_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00010:
        casez_tmp_184 = T_38110_2_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00011:
        casez_tmp_184 = T_38110_3_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00100:
        casez_tmp_184 = T_38110_4_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00101:
        casez_tmp_184 = T_38110_5_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00110:
        casez_tmp_184 = T_38110_6_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b00111:
        casez_tmp_184 = T_38110_7_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01000:
        casez_tmp_184 = T_38110_8_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01001:
        casez_tmp_184 = T_38110_9_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01010:
        casez_tmp_184 = T_38110_10_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01011:
        casez_tmp_184 = T_38110_11_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01100:
        casez_tmp_184 = T_38110_12_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01101:
        casez_tmp_184 = T_38110_13_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01110:
        casez_tmp_184 = T_38110_14_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b01111:
        casez_tmp_184 = T_38110_15_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10000:
        casez_tmp_184 = T_38110_16_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10001:
        casez_tmp_184 = T_38110_17_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10010:
        casez_tmp_184 = T_38110_18_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10011:
        casez_tmp_184 = T_38110_19_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10100:
        casez_tmp_184 = T_38110_20_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10101:
        casez_tmp_184 = T_38110_21_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10110:
        casez_tmp_184 = T_38110_22_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b10111:
        casez_tmp_184 = T_38110_23_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11000:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11001:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11010:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11011:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11100:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11101:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      5'b11110:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
      default:
        casez_tmp_184 = T_38110_0_ldst_val;	// rob.scala:350:34, :531:53, :538:75
    endcase	// rob.scala:531:53, :538:75
  end // always @(*)
  wire _T_47531 = rob_state != 2'h1 & rob_state != 2'h3;	// rob.scala:443:23, :453:100, :574:{34,48,62}, :931:42
  wire _T_3 = _T_29094 & ~_T_29090 & ~_T_47531;	// rob.scala:583:57, :585:{48,72}
  wire _T_47551 = casez_tmp_2 & (~_T_29094 | _T_29090) | _T_47531;	// rob.scala:433:51, :586:48, :587:{31,46,74}
  wire _will_throw_exception = _T_41018 & ~_T_47551 & ~_T_3 | _T_29090 & ~_T_47531;	// rob.scala:514:7, :583:{54,57,71,87}
  wire _T_4 = casez_tmp_94 & ~T_35638_R0_data & ~_T_41018 & ~_T_47551;	// rob.scala:335:30, :433:51, :439:45, :583:57, :585:{48,72}
  wire _T_47568 = _will_throw_exception | io_cxcpt_valid;	// rob.scala:593:48
  wire _T_47569 = r_xcpt_uop_exc_cause == 64'hD;	// rob.scala:594:45, :597:24
  wire [3:0] _rob_head_4to1 = rob_head[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:900:33
  wire _T_47590 = rob_head[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:902:23
  wire _T_5 = _T_47568 | _T_3 & casez_tmp_66 | _T_4 & casez_tmp_158;	// rob.scala:453:59, :608:37, :609:64
  `ifndef SYNTHESIS	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
    `ifdef RANDOMIZE_REG_INIT	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      reg [31:0] _RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      reg [31:0] _RANDOM_233;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_234;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_235;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_236;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_237;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_238;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_239;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_240;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_241;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_242;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_243;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_244;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_245;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_246;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
      reg [31:0] _RANDOM_247;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:38:5
      reg [31:0] _RANDOM_248;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
      reg [31:0] _RANDOM_249;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_250;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_251;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_252;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_253;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_254;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_255;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_256;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_257;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_258;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_259;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_260;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_261;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_262;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_263;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_264;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_265;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_266;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_267;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_268;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_269;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_270;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_271;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_272;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_273;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_274;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_275;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_276;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_277;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_278;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_279;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_280;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_281;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_282;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_283;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_284;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_285;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_286;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_287;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_288;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_289;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_290;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_291;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_292;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_293;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_294;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_295;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_296;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_297;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_298;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_299;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_300;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_301;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_302;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_303;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_304;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_305;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_306;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_307;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_308;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_309;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_310;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_311;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_312;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_313;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_314;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_315;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_316;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_317;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_318;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_319;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_320;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_321;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_322;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_323;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_324;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_325;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_326;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_327;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_328;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_329;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_330;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_331;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_332;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_333;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_334;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_335;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_336;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_337;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_338;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_339;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_340;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_341;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_342;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_343;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_344;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_345;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_346;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_347;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_348;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_349;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_350;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_351;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_352;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_353;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_354;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_355;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_356;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_357;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_358;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_359;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_360;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_361;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_362;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_363;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_364;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_365;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_366;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_367;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_368;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_369;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_370;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_371;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_372;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_373;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_374;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_375;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_376;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_377;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_378;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_379;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_380;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_381;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_382;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_383;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_384;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_385;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_386;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_387;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_388;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_389;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_390;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_391;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_392;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_393;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_394;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_395;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_396;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_397;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_398;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_399;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_400;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_401;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_402;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_403;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_404;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_405;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_406;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_407;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_408;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_409;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_410;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_411;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_412;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_413;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_414;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_415;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_416;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_417;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_418;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_419;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_420;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_421;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_422;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_423;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_424;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_425;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_426;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_427;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_428;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_429;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_430;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_431;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_432;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_433;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_434;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_435;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_436;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_437;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_438;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_439;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_440;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_441;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_442;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_443;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_444;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_445;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_446;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_447;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_448;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_449;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_450;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_451;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_452;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_453;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_454;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_455;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_456;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_457;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_458;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_459;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_460;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_461;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_462;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_463;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_464;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_465;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_466;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_467;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_468;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_469;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_470;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_471;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_472;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_473;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_474;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_475;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_476;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_477;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_478;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_479;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_480;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_481;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_482;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_483;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_484;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_485;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_486;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_487;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_488;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_489;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_490;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_491;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_492;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_493;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_494;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_495;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_496;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_497;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_498;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_499;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_500;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_501;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_502;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_503;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_504;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_505;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_506;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_507;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_508;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_509;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_510;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_511;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_512;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_513;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_514;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_515;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_516;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_517;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_518;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_519;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_520;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_521;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_522;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_523;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_524;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_525;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_526;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_527;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_528;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_529;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_530;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_531;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_532;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_533;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_534;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_535;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_536;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_537;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_538;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_539;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_540;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_541;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_542;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_543;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_544;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_545;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_546;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_547;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_548;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_549;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_550;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_551;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_552;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_553;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_554;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_555;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_556;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_557;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_558;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_559;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_560;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_561;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_562;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_563;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_564;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_565;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_566;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_567;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_568;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_569;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_570;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_571;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_572;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_573;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_574;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_575;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_576;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_577;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_578;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_579;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_580;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_581;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_582;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_583;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_584;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_585;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
      reg [31:0] _RANDOM_586;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_587;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_588;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_589;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_590;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_591;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_592;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_593;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_594;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_595;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_596;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_597;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_598;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_599;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_600;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_601;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_602;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_603;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_604;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_605;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_606;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_607;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_608;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_609;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_610;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_611;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_612;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_613;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_614;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_615;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_616;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_617;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_618;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_619;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_620;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_621;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_622;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_623;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_624;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_625;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_626;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_627;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_628;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_629;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_630;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_631;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_632;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_633;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_634;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_635;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_636;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_637;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_638;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_639;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_640;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_641;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_642;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_643;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_644;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_645;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_646;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_647;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_648;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_649;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_650;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_651;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_652;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_653;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_654;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_655;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_656;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_657;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_658;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_659;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_660;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_661;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_662;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_663;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_664;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_665;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_666;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_667;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_668;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_669;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_670;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_671;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_672;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_673;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_674;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_675;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_676;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_677;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_678;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_679;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_680;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_681;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_682;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_683;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_684;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_685;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_686;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_687;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_688;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_689;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_690;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_691;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_692;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_693;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_694;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_695;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_696;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_697;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_698;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_699;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_700;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_701;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_702;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_703;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_704;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_705;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_706;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_707;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_708;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_709;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_710;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_711;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_712;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_713;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_714;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_715;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_716;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_717;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_718;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_719;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_720;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_721;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_722;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_723;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_724;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_725;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_726;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_727;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_728;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_729;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_730;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_731;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_732;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_733;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_734;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_735;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_736;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_737;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_738;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_739;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_740;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_741;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_742;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_743;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_744;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_745;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_746;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_747;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_748;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_749;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_750;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_751;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_752;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_753;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_754;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_755;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_756;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_757;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_758;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_759;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_760;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_761;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_762;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_763;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_764;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_765;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_766;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_767;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_768;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_769;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_770;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_771;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_772;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_773;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_774;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_775;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_776;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_777;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_778;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_779;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_780;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_781;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_782;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_783;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_784;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_785;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_786;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_787;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_788;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_789;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_790;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_791;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_792;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_793;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_794;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_795;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_796;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_797;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_798;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_799;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_800;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_801;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_802;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_803;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_804;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_805;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_806;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_807;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_808;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_809;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_810;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_811;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_812;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_813;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_814;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_815;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_816;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_817;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_818;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_819;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_820;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_821;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_822;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_823;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_824;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_825;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_826;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_827;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_828;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_829;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_830;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_831;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_832;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_833;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_834;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_835;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_836;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_837;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_838;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_839;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_840;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_841;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_842;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_843;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_844;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_845;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_846;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_847;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_848;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_849;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_850;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_851;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_852;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_853;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_854;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_855;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_856;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_857;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_858;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_859;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_860;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_861;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_862;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_863;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_864;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_865;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_866;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_867;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_868;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_869;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_870;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_871;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_872;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_873;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_874;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_875;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_876;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_877;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_878;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_879;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_880;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_881;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_882;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_883;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_884;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_885;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_886;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_887;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_888;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_889;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_890;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_891;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_892;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_893;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_894;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_895;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_896;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_897;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_898;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_899;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_900;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_901;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_902;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_903;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_904;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_905;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_906;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_907;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_908;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_909;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_910;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_911;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_912;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_913;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_914;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_915;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_916;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_917;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_918;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_919;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_920;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_921;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
      reg [31:0] _RANDOM_922;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5

    `endif
    initial begin	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      `INIT_RANDOM_PROLOG_	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      `ifdef RANDOMIZE_REG_INIT	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
        _RANDOM = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
        rob_state = _RANDOM[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
        rob_head = _RANDOM[6:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:5
        rob_tail = _RANDOM[11:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:14:5
        r_xcpt_val = _RANDOM[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:36:5
        r_xcpt_uop_valid = _RANDOM[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_iw_state = _RANDOM[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_uopc = _RANDOM[24:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_233 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_inst = {_RANDOM_233[24:0], _RANDOM[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_234 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_235 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_pc = {_RANDOM_235[0], _RANDOM_234, _RANDOM_233[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_fu_code = _RANDOM_235[8:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_br_type = _RANDOM_235[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_op1_sel = _RANDOM_235[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_op2_sel = _RANDOM_235[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_imm_sel = _RANDOM_235[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_op_fcn = _RANDOM_235[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_fcn_dw = _RANDOM_235[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_rf_wen = _RANDOM_235[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_csr_cmd = _RANDOM_235[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_is_load = _RANDOM_235[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_is_sta = _RANDOM_235[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_236 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ctrl_is_std = _RANDOM_236[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_wakeup_delay = _RANDOM_236[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_allocate_brtag = _RANDOM_236[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_br_or_jmp = _RANDOM_236[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_jump = _RANDOM_236[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_jal = _RANDOM_236[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_ret = _RANDOM_236[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_call = _RANDOM_236[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_mask = _RANDOM_236[16:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_tag = _RANDOM_236[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_prediction_bpd_predict_val = _RANDOM_236[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_prediction_bpd_predict_taken = _RANDOM_236[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_prediction_btb_hit = _RANDOM_236[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_prediction_btb_predicted = _RANDOM_236[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_br_prediction_is_br_or_jalr = _RANDOM_236[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stat_brjmp_mispredicted = _RANDOM_236[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stat_btb_made_pred = _RANDOM_236[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stat_btb_mispredicted = _RANDOM_236[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stat_bpd_made_pred = _RANDOM_236[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stat_bpd_mispredicted = _RANDOM_236[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_237 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_fetch_pc_lob = {_RANDOM_237[0], _RANDOM_236[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_imm_packed = _RANDOM_237[20:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_238 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_csr_addr = {_RANDOM_238[0], _RANDOM_237[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_rob_idx = _RANDOM_238[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ldq_idx = _RANDOM_238[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stq_idx = _RANDOM_238[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_brob_idx = _RANDOM_238[19:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_pdst = _RANDOM_238[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_239 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_pop1 = {_RANDOM_239[1:0], _RANDOM_238[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_pop2 = _RANDOM_239[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_pop3 = _RANDOM_239[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_prs1_busy = _RANDOM_239[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_prs2_busy = _RANDOM_239[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_prs3_busy = _RANDOM_239[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_stale_pdst = _RANDOM_239[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_exception = _RANDOM_239[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_240 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_241 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_exc_cause = {_RANDOM_241[26:0], _RANDOM_240, _RANDOM_239[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_bypassable = _RANDOM_241[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_mem_cmd = _RANDOM_241[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_242 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_mem_typ = _RANDOM_242[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_fence = _RANDOM_242[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_fencei = _RANDOM_242[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_store = _RANDOM_242[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_amo = _RANDOM_242[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_load = _RANDOM_242[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_is_unique = _RANDOM_242[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_flush_on_commit = _RANDOM_242[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ldst = _RANDOM_242[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_lrs1 = _RANDOM_242[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_lrs2 = _RANDOM_242[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_243 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_lrs3 = {_RANDOM_243[1:0], _RANDOM_242[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_ldst_val = _RANDOM_243[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_dst_rtype = _RANDOM_243[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_lrs1_rtype = _RANDOM_243[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_lrs2_rtype = _RANDOM_243[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_frs3_en = _RANDOM_243[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_fp_val = _RANDOM_243[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_fp_single = _RANDOM_243[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_xcpt_if = _RANDOM_243[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_replay_if = _RANDOM_243[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_244 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_245 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_debug_wdata = {_RANDOM_245[13:0], _RANDOM_244, _RANDOM_243[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_246 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        r_xcpt_uop_debug_events_fetch_seq = {_RANDOM_246[13:0], _RANDOM_245[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:37:5
        _RANDOM_247 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:38:5
        r_xcpt_badvaddr = {_RANDOM_247[21:0], _RANDOM_246[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:38:5
        r_partial_row = _RANDOM_247[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:125:5
        T_23706_0 = _RANDOM_247[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_1 = _RANDOM_247[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_2 = _RANDOM_247[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_3 = _RANDOM_247[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_4 = _RANDOM_247[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_5 = _RANDOM_247[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_6 = _RANDOM_247[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_7 = _RANDOM_247[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_8 = _RANDOM_247[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        _RANDOM_248 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_9 = _RANDOM_248[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_10 = _RANDOM_248[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_11 = _RANDOM_248[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_12 = _RANDOM_248[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_13 = _RANDOM_248[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_14 = _RANDOM_248[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_15 = _RANDOM_248[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_16 = _RANDOM_248[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_17 = _RANDOM_248[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_18 = _RANDOM_248[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_19 = _RANDOM_248[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_20 = _RANDOM_248[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_21 = _RANDOM_248[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_22 = _RANDOM_248[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_23706_23 = _RANDOM_248[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:187:5
        T_26182_0_valid = _RANDOM_248[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_iw_state = _RANDOM_248[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_uopc = _RANDOM_248[26:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_249 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_inst = {_RANDOM_249[26:0], _RANDOM_248[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_250 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_251 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_pc = {_RANDOM_251[2:0], _RANDOM_250, _RANDOM_249[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_fu_code = _RANDOM_251[10:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_br_type = _RANDOM_251[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_op1_sel = _RANDOM_251[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_op2_sel = _RANDOM_251[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_imm_sel = _RANDOM_251[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_op_fcn = _RANDOM_251[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_fcn_dw = _RANDOM_251[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_rf_wen = _RANDOM_251[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_csr_cmd = _RANDOM_251[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_252 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_is_load = _RANDOM_252[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_is_sta = _RANDOM_252[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ctrl_is_std = _RANDOM_252[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_wakeup_delay = _RANDOM_252[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_allocate_brtag = _RANDOM_252[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_br_or_jmp = _RANDOM_252[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_jump = _RANDOM_252[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_jal = _RANDOM_252[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_ret = _RANDOM_252[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_call = _RANDOM_252[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_mask = _RANDOM_252[18:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_tag = _RANDOM_252[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_prediction_bpd_predict_val = _RANDOM_252[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_prediction_bpd_predict_taken = _RANDOM_252[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_prediction_btb_hit = _RANDOM_252[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_prediction_btb_predicted = _RANDOM_252[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_br_prediction_is_br_or_jalr = _RANDOM_252[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stat_brjmp_mispredicted = _RANDOM_252[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stat_btb_made_pred = _RANDOM_252[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stat_btb_mispredicted = _RANDOM_252[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stat_bpd_made_pred = _RANDOM_252[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stat_bpd_mispredicted = _RANDOM_252[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_253 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_fetch_pc_lob = _RANDOM_253[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_imm_packed = _RANDOM_253[22:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_254 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_csr_addr = {_RANDOM_254[2:0], _RANDOM_253[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_rob_idx = _RANDOM_254[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ldq_idx = _RANDOM_254[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stq_idx = _RANDOM_254[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_brob_idx = _RANDOM_254[21:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_pdst = _RANDOM_254[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_255 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_pop1 = {_RANDOM_255[3:0], _RANDOM_254[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_pop2 = _RANDOM_255[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_pop3 = _RANDOM_255[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_prs1_busy = _RANDOM_255[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_prs2_busy = _RANDOM_255[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_prs3_busy = _RANDOM_255[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_stale_pdst = _RANDOM_255[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_exception = _RANDOM_255[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_256 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_257 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_exc_cause = {_RANDOM_257[28:0], _RANDOM_256, _RANDOM_255[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_bypassable = _RANDOM_257[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_258 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_mem_cmd = {_RANDOM_258[1:0], _RANDOM_257[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_mem_typ = _RANDOM_258[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_fence = _RANDOM_258[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_fencei = _RANDOM_258[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_store = _RANDOM_258[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_amo = _RANDOM_258[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_load = _RANDOM_258[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_is_unique = _RANDOM_258[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_flush_on_commit = _RANDOM_258[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ldst = _RANDOM_258[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_lrs1 = _RANDOM_258[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_lrs2 = _RANDOM_258[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_259 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_lrs3 = {_RANDOM_259[3:0], _RANDOM_258[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_ldst_val = _RANDOM_259[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_dst_rtype = _RANDOM_259[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_lrs1_rtype = _RANDOM_259[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_lrs2_rtype = _RANDOM_259[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_frs3_en = _RANDOM_259[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_fp_val = _RANDOM_259[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_fp_single = _RANDOM_259[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_xcpt_if = _RANDOM_259[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_replay_if = _RANDOM_259[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_260 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_261 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_debug_wdata = {_RANDOM_261[15:0], _RANDOM_260, _RANDOM_259[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_262 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_0_debug_events_fetch_seq = {_RANDOM_262[15:0], _RANDOM_261[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_valid = _RANDOM_262[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_iw_state = _RANDOM_262[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_uopc = _RANDOM_262[27:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_263 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_inst = {_RANDOM_263[27:0], _RANDOM_262[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_264 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_265 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_pc = {_RANDOM_265[3:0], _RANDOM_264, _RANDOM_263[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_fu_code = _RANDOM_265[11:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_br_type = _RANDOM_265[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_op1_sel = _RANDOM_265[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_op2_sel = _RANDOM_265[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_imm_sel = _RANDOM_265[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_op_fcn = _RANDOM_265[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_fcn_dw = _RANDOM_265[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_rf_wen = _RANDOM_265[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_266 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_csr_cmd = {_RANDOM_266[0], _RANDOM_265[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_is_load = _RANDOM_266[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_is_sta = _RANDOM_266[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ctrl_is_std = _RANDOM_266[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_wakeup_delay = _RANDOM_266[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_allocate_brtag = _RANDOM_266[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_br_or_jmp = _RANDOM_266[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_jump = _RANDOM_266[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_jal = _RANDOM_266[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_ret = _RANDOM_266[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_call = _RANDOM_266[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_mask = _RANDOM_266[19:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_tag = _RANDOM_266[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_prediction_bpd_predict_val = _RANDOM_266[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_prediction_bpd_predict_taken = _RANDOM_266[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_prediction_btb_hit = _RANDOM_266[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_prediction_btb_predicted = _RANDOM_266[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_br_prediction_is_br_or_jalr = _RANDOM_266[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stat_brjmp_mispredicted = _RANDOM_266[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stat_btb_made_pred = _RANDOM_266[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stat_btb_mispredicted = _RANDOM_266[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stat_bpd_made_pred = _RANDOM_266[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_267 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stat_bpd_mispredicted = _RANDOM_267[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_fetch_pc_lob = _RANDOM_267[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_imm_packed = _RANDOM_267[23:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_268 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_csr_addr = {_RANDOM_268[3:0], _RANDOM_267[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_rob_idx = _RANDOM_268[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ldq_idx = _RANDOM_268[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stq_idx = _RANDOM_268[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_brob_idx = _RANDOM_268[22:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_pdst = _RANDOM_268[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_269 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_pop1 = {_RANDOM_269[4:0], _RANDOM_268[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_pop2 = _RANDOM_269[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_pop3 = _RANDOM_269[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_prs1_busy = _RANDOM_269[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_prs2_busy = _RANDOM_269[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_prs3_busy = _RANDOM_269[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_stale_pdst = _RANDOM_269[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_exception = _RANDOM_269[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_270 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_271 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_exc_cause = {_RANDOM_271[29:0], _RANDOM_270, _RANDOM_269[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_bypassable = _RANDOM_271[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_272 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_mem_cmd = {_RANDOM_272[2:0], _RANDOM_271[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_mem_typ = _RANDOM_272[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_fence = _RANDOM_272[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_fencei = _RANDOM_272[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_store = _RANDOM_272[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_amo = _RANDOM_272[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_load = _RANDOM_272[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_is_unique = _RANDOM_272[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_flush_on_commit = _RANDOM_272[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ldst = _RANDOM_272[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_lrs1 = _RANDOM_272[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_lrs2 = _RANDOM_272[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_273 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_lrs3 = {_RANDOM_273[4:0], _RANDOM_272[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_ldst_val = _RANDOM_273[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_dst_rtype = _RANDOM_273[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_lrs1_rtype = _RANDOM_273[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_lrs2_rtype = _RANDOM_273[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_frs3_en = _RANDOM_273[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_fp_val = _RANDOM_273[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_fp_single = _RANDOM_273[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_xcpt_if = _RANDOM_273[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_replay_if = _RANDOM_273[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_274 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_275 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_debug_wdata = {_RANDOM_275[16:0], _RANDOM_274, _RANDOM_273[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_276 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_1_debug_events_fetch_seq = {_RANDOM_276[16:0], _RANDOM_275[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_valid = _RANDOM_276[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_iw_state = _RANDOM_276[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_uopc = _RANDOM_276[28:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_277 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_inst = {_RANDOM_277[28:0], _RANDOM_276[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_278 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_279 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_pc = {_RANDOM_279[4:0], _RANDOM_278, _RANDOM_277[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_fu_code = _RANDOM_279[12:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_br_type = _RANDOM_279[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_op1_sel = _RANDOM_279[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_op2_sel = _RANDOM_279[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_imm_sel = _RANDOM_279[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_op_fcn = _RANDOM_279[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_fcn_dw = _RANDOM_279[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_rf_wen = _RANDOM_279[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_280 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_csr_cmd = {_RANDOM_280[1:0], _RANDOM_279[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_is_load = _RANDOM_280[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_is_sta = _RANDOM_280[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ctrl_is_std = _RANDOM_280[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_wakeup_delay = _RANDOM_280[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_allocate_brtag = _RANDOM_280[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_br_or_jmp = _RANDOM_280[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_jump = _RANDOM_280[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_jal = _RANDOM_280[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_ret = _RANDOM_280[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_call = _RANDOM_280[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_mask = _RANDOM_280[20:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_tag = _RANDOM_280[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_prediction_bpd_predict_val = _RANDOM_280[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_prediction_bpd_predict_taken = _RANDOM_280[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_prediction_btb_hit = _RANDOM_280[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_prediction_btb_predicted = _RANDOM_280[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_br_prediction_is_br_or_jalr = _RANDOM_280[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stat_brjmp_mispredicted = _RANDOM_280[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stat_btb_made_pred = _RANDOM_280[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stat_btb_mispredicted = _RANDOM_280[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_281 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stat_bpd_made_pred = _RANDOM_281[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stat_bpd_mispredicted = _RANDOM_281[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_fetch_pc_lob = _RANDOM_281[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_imm_packed = _RANDOM_281[24:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_282 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_csr_addr = {_RANDOM_282[4:0], _RANDOM_281[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_rob_idx = _RANDOM_282[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ldq_idx = _RANDOM_282[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stq_idx = _RANDOM_282[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_brob_idx = _RANDOM_282[23:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_pdst = _RANDOM_282[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_283 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_pop1 = {_RANDOM_283[5:0], _RANDOM_282[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_pop2 = _RANDOM_283[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_pop3 = _RANDOM_283[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_prs1_busy = _RANDOM_283[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_prs2_busy = _RANDOM_283[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_prs3_busy = _RANDOM_283[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_stale_pdst = _RANDOM_283[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_exception = _RANDOM_283[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_284 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_285 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_exc_cause = {_RANDOM_285[30:0], _RANDOM_284, _RANDOM_283[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_bypassable = _RANDOM_285[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_286 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_mem_cmd = _RANDOM_286[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_mem_typ = _RANDOM_286[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_fence = _RANDOM_286[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_fencei = _RANDOM_286[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_store = _RANDOM_286[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_amo = _RANDOM_286[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_load = _RANDOM_286[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_is_unique = _RANDOM_286[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_flush_on_commit = _RANDOM_286[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ldst = _RANDOM_286[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_lrs1 = _RANDOM_286[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_lrs2 = _RANDOM_286[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_287 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_lrs3 = _RANDOM_287[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_ldst_val = _RANDOM_287[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_dst_rtype = _RANDOM_287[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_lrs1_rtype = _RANDOM_287[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_lrs2_rtype = _RANDOM_287[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_frs3_en = _RANDOM_287[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_fp_val = _RANDOM_287[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_fp_single = _RANDOM_287[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_xcpt_if = _RANDOM_287[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_replay_if = _RANDOM_287[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_288 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_289 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_debug_wdata = {_RANDOM_289[17:0], _RANDOM_288, _RANDOM_287[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_290 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_2_debug_events_fetch_seq = {_RANDOM_290[17:0], _RANDOM_289[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_valid = _RANDOM_290[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_iw_state = _RANDOM_290[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_uopc = _RANDOM_290[29:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_291 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_inst = {_RANDOM_291[29:0], _RANDOM_290[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_292 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_293 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_pc = {_RANDOM_293[5:0], _RANDOM_292, _RANDOM_291[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_fu_code = _RANDOM_293[13:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_br_type = _RANDOM_293[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_op1_sel = _RANDOM_293[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_op2_sel = _RANDOM_293[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_imm_sel = _RANDOM_293[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_op_fcn = _RANDOM_293[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_fcn_dw = _RANDOM_293[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_rf_wen = _RANDOM_293[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_294 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_csr_cmd = _RANDOM_294[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_is_load = _RANDOM_294[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_is_sta = _RANDOM_294[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ctrl_is_std = _RANDOM_294[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_wakeup_delay = _RANDOM_294[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_allocate_brtag = _RANDOM_294[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_br_or_jmp = _RANDOM_294[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_jump = _RANDOM_294[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_jal = _RANDOM_294[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_ret = _RANDOM_294[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_call = _RANDOM_294[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_mask = _RANDOM_294[21:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_tag = _RANDOM_294[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_prediction_bpd_predict_val = _RANDOM_294[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_prediction_bpd_predict_taken = _RANDOM_294[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_prediction_btb_hit = _RANDOM_294[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_prediction_btb_predicted = _RANDOM_294[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_br_prediction_is_br_or_jalr = _RANDOM_294[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stat_brjmp_mispredicted = _RANDOM_294[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stat_btb_made_pred = _RANDOM_294[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_295 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stat_btb_mispredicted = _RANDOM_295[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stat_bpd_made_pred = _RANDOM_295[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stat_bpd_mispredicted = _RANDOM_295[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_fetch_pc_lob = _RANDOM_295[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_imm_packed = _RANDOM_295[25:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_296 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_csr_addr = {_RANDOM_296[5:0], _RANDOM_295[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_rob_idx = _RANDOM_296[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ldq_idx = _RANDOM_296[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stq_idx = _RANDOM_296[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_brob_idx = _RANDOM_296[24:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_pdst = _RANDOM_296[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_297 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_pop1 = _RANDOM_297[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_pop2 = _RANDOM_297[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_pop3 = _RANDOM_297[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_prs1_busy = _RANDOM_297[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_prs2_busy = _RANDOM_297[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_prs3_busy = _RANDOM_297[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_stale_pdst = _RANDOM_297[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_exception = _RANDOM_297[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_298 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_299 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_exc_cause = {_RANDOM_299, _RANDOM_298};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_300 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_bypassable = _RANDOM_300[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_mem_cmd = _RANDOM_300[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_mem_typ = _RANDOM_300[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_fence = _RANDOM_300[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_fencei = _RANDOM_300[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_store = _RANDOM_300[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_amo = _RANDOM_300[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_load = _RANDOM_300[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_is_unique = _RANDOM_300[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_flush_on_commit = _RANDOM_300[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ldst = _RANDOM_300[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_lrs1 = _RANDOM_300[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_301 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_lrs2 = {_RANDOM_301[0], _RANDOM_300[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_lrs3 = _RANDOM_301[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_ldst_val = _RANDOM_301[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_dst_rtype = _RANDOM_301[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_lrs1_rtype = _RANDOM_301[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_lrs2_rtype = _RANDOM_301[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_frs3_en = _RANDOM_301[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_fp_val = _RANDOM_301[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_fp_single = _RANDOM_301[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_xcpt_if = _RANDOM_301[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_replay_if = _RANDOM_301[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_302 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_303 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_debug_wdata = {_RANDOM_303[18:0], _RANDOM_302, _RANDOM_301[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_304 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_3_debug_events_fetch_seq = {_RANDOM_304[18:0], _RANDOM_303[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_valid = _RANDOM_304[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_iw_state = _RANDOM_304[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_uopc = _RANDOM_304[30:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_305 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_inst = {_RANDOM_305[30:0], _RANDOM_304[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_306 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_307 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_pc = {_RANDOM_307[6:0], _RANDOM_306, _RANDOM_305[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_fu_code = _RANDOM_307[14:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_br_type = _RANDOM_307[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_op1_sel = _RANDOM_307[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_op2_sel = _RANDOM_307[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_imm_sel = _RANDOM_307[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_op_fcn = _RANDOM_307[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_fcn_dw = _RANDOM_307[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_308 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_rf_wen = _RANDOM_308[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_csr_cmd = _RANDOM_308[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_is_load = _RANDOM_308[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_is_sta = _RANDOM_308[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ctrl_is_std = _RANDOM_308[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_wakeup_delay = _RANDOM_308[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_allocate_brtag = _RANDOM_308[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_br_or_jmp = _RANDOM_308[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_jump = _RANDOM_308[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_jal = _RANDOM_308[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_ret = _RANDOM_308[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_call = _RANDOM_308[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_mask = _RANDOM_308[22:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_tag = _RANDOM_308[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_prediction_bpd_predict_val = _RANDOM_308[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_prediction_bpd_predict_taken = _RANDOM_308[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_prediction_btb_hit = _RANDOM_308[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_prediction_btb_predicted = _RANDOM_308[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_br_prediction_is_br_or_jalr = _RANDOM_308[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stat_brjmp_mispredicted = _RANDOM_308[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_309 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stat_btb_made_pred = _RANDOM_309[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stat_btb_mispredicted = _RANDOM_309[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stat_bpd_made_pred = _RANDOM_309[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stat_bpd_mispredicted = _RANDOM_309[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_fetch_pc_lob = _RANDOM_309[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_imm_packed = _RANDOM_309[26:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_310 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_csr_addr = {_RANDOM_310[6:0], _RANDOM_309[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_rob_idx = _RANDOM_310[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ldq_idx = _RANDOM_310[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stq_idx = _RANDOM_310[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_brob_idx = _RANDOM_310[25:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_311 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_pdst = {_RANDOM_311[0], _RANDOM_310[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_pop1 = _RANDOM_311[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_pop2 = _RANDOM_311[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_pop3 = _RANDOM_311[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_prs1_busy = _RANDOM_311[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_prs2_busy = _RANDOM_311[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_prs3_busy = _RANDOM_311[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_stale_pdst = _RANDOM_311[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_312 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_exception = _RANDOM_312[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_313 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_314 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_exc_cause = {_RANDOM_314[0], _RANDOM_313, _RANDOM_312[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_bypassable = _RANDOM_314[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_mem_cmd = _RANDOM_314[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_mem_typ = _RANDOM_314[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_fence = _RANDOM_314[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_fencei = _RANDOM_314[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_store = _RANDOM_314[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_amo = _RANDOM_314[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_load = _RANDOM_314[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_is_unique = _RANDOM_314[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_flush_on_commit = _RANDOM_314[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ldst = _RANDOM_314[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_lrs1 = _RANDOM_314[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_315 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_lrs2 = {_RANDOM_315[1:0], _RANDOM_314[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_lrs3 = _RANDOM_315[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_ldst_val = _RANDOM_315[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_dst_rtype = _RANDOM_315[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_lrs1_rtype = _RANDOM_315[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_lrs2_rtype = _RANDOM_315[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_frs3_en = _RANDOM_315[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_fp_val = _RANDOM_315[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_fp_single = _RANDOM_315[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_xcpt_if = _RANDOM_315[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_replay_if = _RANDOM_315[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_316 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_317 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_debug_wdata = {_RANDOM_317[19:0], _RANDOM_316, _RANDOM_315[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_318 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_4_debug_events_fetch_seq = {_RANDOM_318[19:0], _RANDOM_317[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_valid = _RANDOM_318[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_iw_state = _RANDOM_318[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_uopc = _RANDOM_318[31:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_319 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_inst = _RANDOM_319;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_320 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_321 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_pc = {_RANDOM_321[7:0], _RANDOM_320};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_fu_code = _RANDOM_321[15:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_br_type = _RANDOM_321[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_op1_sel = _RANDOM_321[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_op2_sel = _RANDOM_321[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_imm_sel = _RANDOM_321[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_op_fcn = _RANDOM_321[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_322 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_fcn_dw = _RANDOM_322[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_rf_wen = _RANDOM_322[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_csr_cmd = _RANDOM_322[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_is_load = _RANDOM_322[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_is_sta = _RANDOM_322[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ctrl_is_std = _RANDOM_322[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_wakeup_delay = _RANDOM_322[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_allocate_brtag = _RANDOM_322[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_br_or_jmp = _RANDOM_322[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_jump = _RANDOM_322[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_jal = _RANDOM_322[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_ret = _RANDOM_322[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_call = _RANDOM_322[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_mask = _RANDOM_322[23:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_tag = _RANDOM_322[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_prediction_bpd_predict_val = _RANDOM_322[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_prediction_bpd_predict_taken = _RANDOM_322[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_prediction_btb_hit = _RANDOM_322[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_prediction_btb_predicted = _RANDOM_322[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_br_prediction_is_br_or_jalr = _RANDOM_322[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_323 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stat_brjmp_mispredicted = _RANDOM_323[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stat_btb_made_pred = _RANDOM_323[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stat_btb_mispredicted = _RANDOM_323[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stat_bpd_made_pred = _RANDOM_323[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stat_bpd_mispredicted = _RANDOM_323[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_fetch_pc_lob = _RANDOM_323[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_imm_packed = _RANDOM_323[27:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_324 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_csr_addr = {_RANDOM_324[7:0], _RANDOM_323[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_rob_idx = _RANDOM_324[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ldq_idx = _RANDOM_324[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stq_idx = _RANDOM_324[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_brob_idx = _RANDOM_324[26:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_325 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_pdst = {_RANDOM_325[1:0], _RANDOM_324[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_pop1 = _RANDOM_325[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_pop2 = _RANDOM_325[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_pop3 = _RANDOM_325[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_prs1_busy = _RANDOM_325[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_prs2_busy = _RANDOM_325[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_prs3_busy = _RANDOM_325[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_326 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_stale_pdst = {_RANDOM_326[0], _RANDOM_325[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_exception = _RANDOM_326[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_327 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_328 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_exc_cause = {_RANDOM_328[1:0], _RANDOM_327, _RANDOM_326[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_bypassable = _RANDOM_328[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_mem_cmd = _RANDOM_328[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_mem_typ = _RANDOM_328[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_fence = _RANDOM_328[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_fencei = _RANDOM_328[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_store = _RANDOM_328[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_amo = _RANDOM_328[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_load = _RANDOM_328[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_is_unique = _RANDOM_328[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_flush_on_commit = _RANDOM_328[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ldst = _RANDOM_328[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_lrs1 = _RANDOM_328[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_329 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_lrs2 = {_RANDOM_329[2:0], _RANDOM_328[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_lrs3 = _RANDOM_329[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_ldst_val = _RANDOM_329[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_dst_rtype = _RANDOM_329[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_lrs1_rtype = _RANDOM_329[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_lrs2_rtype = _RANDOM_329[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_frs3_en = _RANDOM_329[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_fp_val = _RANDOM_329[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_fp_single = _RANDOM_329[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_xcpt_if = _RANDOM_329[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_replay_if = _RANDOM_329[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_330 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_331 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_debug_wdata = {_RANDOM_331[20:0], _RANDOM_330, _RANDOM_329[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_332 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_5_debug_events_fetch_seq = {_RANDOM_332[20:0], _RANDOM_331[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_valid = _RANDOM_332[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_iw_state = _RANDOM_332[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_333 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_uopc = {_RANDOM_333[0], _RANDOM_332[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_334 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_inst = {_RANDOM_334[0], _RANDOM_333[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_335 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_pc = {_RANDOM_335[8:0], _RANDOM_334[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_fu_code = _RANDOM_335[16:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_br_type = _RANDOM_335[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_op1_sel = _RANDOM_335[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_op2_sel = _RANDOM_335[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_imm_sel = _RANDOM_335[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_336 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_op_fcn = {_RANDOM_336[0], _RANDOM_335[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_fcn_dw = _RANDOM_336[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_rf_wen = _RANDOM_336[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_csr_cmd = _RANDOM_336[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_is_load = _RANDOM_336[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_is_sta = _RANDOM_336[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ctrl_is_std = _RANDOM_336[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_wakeup_delay = _RANDOM_336[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_allocate_brtag = _RANDOM_336[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_br_or_jmp = _RANDOM_336[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_jump = _RANDOM_336[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_jal = _RANDOM_336[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_ret = _RANDOM_336[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_call = _RANDOM_336[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_mask = _RANDOM_336[24:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_tag = _RANDOM_336[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_prediction_bpd_predict_val = _RANDOM_336[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_prediction_bpd_predict_taken = _RANDOM_336[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_prediction_btb_hit = _RANDOM_336[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_prediction_btb_predicted = _RANDOM_336[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_337 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_br_prediction_is_br_or_jalr = _RANDOM_337[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stat_brjmp_mispredicted = _RANDOM_337[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stat_btb_made_pred = _RANDOM_337[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stat_btb_mispredicted = _RANDOM_337[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stat_bpd_made_pred = _RANDOM_337[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stat_bpd_mispredicted = _RANDOM_337[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_fetch_pc_lob = _RANDOM_337[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_imm_packed = _RANDOM_337[28:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_338 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_csr_addr = {_RANDOM_338[8:0], _RANDOM_337[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_rob_idx = _RANDOM_338[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ldq_idx = _RANDOM_338[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stq_idx = _RANDOM_338[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_brob_idx = _RANDOM_338[27:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_339 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_pdst = {_RANDOM_339[2:0], _RANDOM_338[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_pop1 = _RANDOM_339[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_pop2 = _RANDOM_339[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_pop3 = _RANDOM_339[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_prs1_busy = _RANDOM_339[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_prs2_busy = _RANDOM_339[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_prs3_busy = _RANDOM_339[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_340 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_stale_pdst = {_RANDOM_340[1:0], _RANDOM_339[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_exception = _RANDOM_340[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_341 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_342 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_exc_cause = {_RANDOM_342[2:0], _RANDOM_341, _RANDOM_340[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_bypassable = _RANDOM_342[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_mem_cmd = _RANDOM_342[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_mem_typ = _RANDOM_342[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_fence = _RANDOM_342[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_fencei = _RANDOM_342[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_store = _RANDOM_342[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_amo = _RANDOM_342[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_load = _RANDOM_342[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_is_unique = _RANDOM_342[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_flush_on_commit = _RANDOM_342[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ldst = _RANDOM_342[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_lrs1 = _RANDOM_342[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_343 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_lrs2 = {_RANDOM_343[3:0], _RANDOM_342[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_lrs3 = _RANDOM_343[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_ldst_val = _RANDOM_343[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_dst_rtype = _RANDOM_343[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_lrs1_rtype = _RANDOM_343[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_lrs2_rtype = _RANDOM_343[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_frs3_en = _RANDOM_343[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_fp_val = _RANDOM_343[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_fp_single = _RANDOM_343[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_xcpt_if = _RANDOM_343[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_replay_if = _RANDOM_343[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_344 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_345 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_debug_wdata = {_RANDOM_345[21:0], _RANDOM_344, _RANDOM_343[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_346 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_6_debug_events_fetch_seq = {_RANDOM_346[21:0], _RANDOM_345[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_valid = _RANDOM_346[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_iw_state = _RANDOM_346[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_347 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_uopc = {_RANDOM_347[1:0], _RANDOM_346[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_348 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_inst = {_RANDOM_348[1:0], _RANDOM_347[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_349 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_pc = {_RANDOM_349[9:0], _RANDOM_348[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_fu_code = _RANDOM_349[17:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_br_type = _RANDOM_349[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_op1_sel = _RANDOM_349[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_op2_sel = _RANDOM_349[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_imm_sel = _RANDOM_349[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_350 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_op_fcn = {_RANDOM_350[1:0], _RANDOM_349[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_fcn_dw = _RANDOM_350[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_rf_wen = _RANDOM_350[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_csr_cmd = _RANDOM_350[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_is_load = _RANDOM_350[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_is_sta = _RANDOM_350[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ctrl_is_std = _RANDOM_350[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_wakeup_delay = _RANDOM_350[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_allocate_brtag = _RANDOM_350[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_br_or_jmp = _RANDOM_350[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_jump = _RANDOM_350[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_jal = _RANDOM_350[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_ret = _RANDOM_350[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_call = _RANDOM_350[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_mask = _RANDOM_350[25:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_tag = _RANDOM_350[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_prediction_bpd_predict_val = _RANDOM_350[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_prediction_bpd_predict_taken = _RANDOM_350[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_prediction_btb_hit = _RANDOM_350[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_351 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_prediction_btb_predicted = _RANDOM_351[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_br_prediction_is_br_or_jalr = _RANDOM_351[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stat_brjmp_mispredicted = _RANDOM_351[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stat_btb_made_pred = _RANDOM_351[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stat_btb_mispredicted = _RANDOM_351[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stat_bpd_made_pred = _RANDOM_351[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stat_bpd_mispredicted = _RANDOM_351[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_fetch_pc_lob = _RANDOM_351[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_imm_packed = _RANDOM_351[29:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_352 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_csr_addr = {_RANDOM_352[9:0], _RANDOM_351[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_rob_idx = _RANDOM_352[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ldq_idx = _RANDOM_352[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stq_idx = _RANDOM_352[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_brob_idx = _RANDOM_352[28:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_353 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_pdst = {_RANDOM_353[3:0], _RANDOM_352[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_pop1 = _RANDOM_353[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_pop2 = _RANDOM_353[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_pop3 = _RANDOM_353[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_prs1_busy = _RANDOM_353[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_prs2_busy = _RANDOM_353[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_prs3_busy = _RANDOM_353[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_354 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_stale_pdst = {_RANDOM_354[2:0], _RANDOM_353[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_exception = _RANDOM_354[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_355 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_356 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_exc_cause = {_RANDOM_356[3:0], _RANDOM_355, _RANDOM_354[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_bypassable = _RANDOM_356[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_mem_cmd = _RANDOM_356[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_mem_typ = _RANDOM_356[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_fence = _RANDOM_356[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_fencei = _RANDOM_356[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_store = _RANDOM_356[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_amo = _RANDOM_356[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_load = _RANDOM_356[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_is_unique = _RANDOM_356[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_flush_on_commit = _RANDOM_356[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ldst = _RANDOM_356[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_lrs1 = _RANDOM_356[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_357 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_lrs2 = {_RANDOM_357[4:0], _RANDOM_356[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_lrs3 = _RANDOM_357[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_ldst_val = _RANDOM_357[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_dst_rtype = _RANDOM_357[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_lrs1_rtype = _RANDOM_357[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_lrs2_rtype = _RANDOM_357[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_frs3_en = _RANDOM_357[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_fp_val = _RANDOM_357[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_fp_single = _RANDOM_357[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_xcpt_if = _RANDOM_357[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_replay_if = _RANDOM_357[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_358 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_359 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_debug_wdata = {_RANDOM_359[22:0], _RANDOM_358, _RANDOM_357[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_360 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_7_debug_events_fetch_seq = {_RANDOM_360[22:0], _RANDOM_359[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_valid = _RANDOM_360[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_iw_state = _RANDOM_360[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_361 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_uopc = {_RANDOM_361[2:0], _RANDOM_360[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_362 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_inst = {_RANDOM_362[2:0], _RANDOM_361[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_363 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_pc = {_RANDOM_363[10:0], _RANDOM_362[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_fu_code = _RANDOM_363[18:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_br_type = _RANDOM_363[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_op1_sel = _RANDOM_363[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_op2_sel = _RANDOM_363[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_imm_sel = _RANDOM_363[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_364 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_op_fcn = {_RANDOM_364[2:0], _RANDOM_363[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_fcn_dw = _RANDOM_364[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_rf_wen = _RANDOM_364[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_csr_cmd = _RANDOM_364[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_is_load = _RANDOM_364[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_is_sta = _RANDOM_364[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ctrl_is_std = _RANDOM_364[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_wakeup_delay = _RANDOM_364[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_allocate_brtag = _RANDOM_364[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_br_or_jmp = _RANDOM_364[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_jump = _RANDOM_364[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_jal = _RANDOM_364[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_ret = _RANDOM_364[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_call = _RANDOM_364[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_mask = _RANDOM_364[26:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_tag = _RANDOM_364[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_prediction_bpd_predict_val = _RANDOM_364[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_prediction_bpd_predict_taken = _RANDOM_364[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_365 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_prediction_btb_hit = _RANDOM_365[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_prediction_btb_predicted = _RANDOM_365[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_br_prediction_is_br_or_jalr = _RANDOM_365[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stat_brjmp_mispredicted = _RANDOM_365[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stat_btb_made_pred = _RANDOM_365[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stat_btb_mispredicted = _RANDOM_365[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stat_bpd_made_pred = _RANDOM_365[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stat_bpd_mispredicted = _RANDOM_365[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_fetch_pc_lob = _RANDOM_365[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_imm_packed = _RANDOM_365[30:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_366 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_csr_addr = {_RANDOM_366[10:0], _RANDOM_365[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_rob_idx = _RANDOM_366[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ldq_idx = _RANDOM_366[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stq_idx = _RANDOM_366[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_brob_idx = _RANDOM_366[29:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_367 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_pdst = {_RANDOM_367[4:0], _RANDOM_366[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_pop1 = _RANDOM_367[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_pop2 = _RANDOM_367[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_pop3 = _RANDOM_367[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_prs1_busy = _RANDOM_367[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_prs2_busy = _RANDOM_367[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_prs3_busy = _RANDOM_367[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_368 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_stale_pdst = {_RANDOM_368[3:0], _RANDOM_367[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_exception = _RANDOM_368[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_369 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_370 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_exc_cause = {_RANDOM_370[4:0], _RANDOM_369, _RANDOM_368[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_bypassable = _RANDOM_370[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_mem_cmd = _RANDOM_370[9:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_mem_typ = _RANDOM_370[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_fence = _RANDOM_370[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_fencei = _RANDOM_370[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_store = _RANDOM_370[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_amo = _RANDOM_370[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_load = _RANDOM_370[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_is_unique = _RANDOM_370[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_flush_on_commit = _RANDOM_370[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ldst = _RANDOM_370[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_lrs1 = _RANDOM_370[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_371 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_lrs2 = _RANDOM_371[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_lrs3 = _RANDOM_371[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_ldst_val = _RANDOM_371[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_dst_rtype = _RANDOM_371[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_lrs1_rtype = _RANDOM_371[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_lrs2_rtype = _RANDOM_371[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_frs3_en = _RANDOM_371[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_fp_val = _RANDOM_371[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_fp_single = _RANDOM_371[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_xcpt_if = _RANDOM_371[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_replay_if = _RANDOM_371[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_372 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_373 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_debug_wdata = {_RANDOM_373[23:0], _RANDOM_372, _RANDOM_371[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_374 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_8_debug_events_fetch_seq = {_RANDOM_374[23:0], _RANDOM_373[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_valid = _RANDOM_374[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_iw_state = _RANDOM_374[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_375 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_uopc = {_RANDOM_375[3:0], _RANDOM_374[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_376 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_inst = {_RANDOM_376[3:0], _RANDOM_375[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_377 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_pc = {_RANDOM_377[11:0], _RANDOM_376[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_fu_code = _RANDOM_377[19:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_br_type = _RANDOM_377[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_op1_sel = _RANDOM_377[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_op2_sel = _RANDOM_377[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_imm_sel = _RANDOM_377[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_378 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_op_fcn = _RANDOM_378[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_fcn_dw = _RANDOM_378[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_rf_wen = _RANDOM_378[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_csr_cmd = _RANDOM_378[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_is_load = _RANDOM_378[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_is_sta = _RANDOM_378[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ctrl_is_std = _RANDOM_378[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_wakeup_delay = _RANDOM_378[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_allocate_brtag = _RANDOM_378[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_br_or_jmp = _RANDOM_378[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_jump = _RANDOM_378[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_jal = _RANDOM_378[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_ret = _RANDOM_378[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_call = _RANDOM_378[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_mask = _RANDOM_378[27:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_tag = _RANDOM_378[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_prediction_bpd_predict_val = _RANDOM_378[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_379 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_prediction_bpd_predict_taken = _RANDOM_379[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_prediction_btb_hit = _RANDOM_379[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_prediction_btb_predicted = _RANDOM_379[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_br_prediction_is_br_or_jalr = _RANDOM_379[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stat_brjmp_mispredicted = _RANDOM_379[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stat_btb_made_pred = _RANDOM_379[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stat_btb_mispredicted = _RANDOM_379[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stat_bpd_made_pred = _RANDOM_379[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stat_bpd_mispredicted = _RANDOM_379[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_fetch_pc_lob = _RANDOM_379[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_imm_packed = _RANDOM_379[31:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_380 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_csr_addr = _RANDOM_380[11:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_rob_idx = _RANDOM_380[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ldq_idx = _RANDOM_380[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stq_idx = _RANDOM_380[25:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_brob_idx = _RANDOM_380[30:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_381 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_pdst = {_RANDOM_381[5:0], _RANDOM_380[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_pop1 = _RANDOM_381[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_pop2 = _RANDOM_381[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_pop3 = _RANDOM_381[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_prs1_busy = _RANDOM_381[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_prs2_busy = _RANDOM_381[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_prs3_busy = _RANDOM_381[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_382 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_stale_pdst = {_RANDOM_382[4:0], _RANDOM_381[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_exception = _RANDOM_382[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_383 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_384 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_exc_cause = {_RANDOM_384[5:0], _RANDOM_383, _RANDOM_382[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_bypassable = _RANDOM_384[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_mem_cmd = _RANDOM_384[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_mem_typ = _RANDOM_384[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_fence = _RANDOM_384[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_fencei = _RANDOM_384[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_store = _RANDOM_384[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_amo = _RANDOM_384[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_load = _RANDOM_384[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_is_unique = _RANDOM_384[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_flush_on_commit = _RANDOM_384[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ldst = _RANDOM_384[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_385 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_lrs1 = {_RANDOM_385[0], _RANDOM_384[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_lrs2 = _RANDOM_385[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_lrs3 = _RANDOM_385[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_ldst_val = _RANDOM_385[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_dst_rtype = _RANDOM_385[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_lrs1_rtype = _RANDOM_385[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_lrs2_rtype = _RANDOM_385[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_frs3_en = _RANDOM_385[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_fp_val = _RANDOM_385[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_fp_single = _RANDOM_385[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_xcpt_if = _RANDOM_385[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_replay_if = _RANDOM_385[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_386 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_387 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_debug_wdata = {_RANDOM_387[24:0], _RANDOM_386, _RANDOM_385[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_388 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_9_debug_events_fetch_seq = {_RANDOM_388[24:0], _RANDOM_387[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_valid = _RANDOM_388[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_iw_state = _RANDOM_388[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_389 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_uopc = {_RANDOM_389[4:0], _RANDOM_388[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_390 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_inst = {_RANDOM_390[4:0], _RANDOM_389[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_391 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_pc = {_RANDOM_391[12:0], _RANDOM_390[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_fu_code = _RANDOM_391[20:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_br_type = _RANDOM_391[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_op1_sel = _RANDOM_391[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_op2_sel = _RANDOM_391[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_392 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_imm_sel = {_RANDOM_392[0], _RANDOM_391[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_op_fcn = _RANDOM_392[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_fcn_dw = _RANDOM_392[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_rf_wen = _RANDOM_392[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_csr_cmd = _RANDOM_392[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_is_load = _RANDOM_392[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_is_sta = _RANDOM_392[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ctrl_is_std = _RANDOM_392[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_wakeup_delay = _RANDOM_392[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_allocate_brtag = _RANDOM_392[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_br_or_jmp = _RANDOM_392[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_jump = _RANDOM_392[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_jal = _RANDOM_392[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_ret = _RANDOM_392[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_call = _RANDOM_392[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_mask = _RANDOM_392[28:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_tag = _RANDOM_392[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_393 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_prediction_bpd_predict_val = _RANDOM_393[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_prediction_bpd_predict_taken = _RANDOM_393[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_prediction_btb_hit = _RANDOM_393[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_prediction_btb_predicted = _RANDOM_393[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_br_prediction_is_br_or_jalr = _RANDOM_393[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stat_brjmp_mispredicted = _RANDOM_393[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stat_btb_made_pred = _RANDOM_393[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stat_btb_mispredicted = _RANDOM_393[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stat_bpd_made_pred = _RANDOM_393[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stat_bpd_mispredicted = _RANDOM_393[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_fetch_pc_lob = _RANDOM_393[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_394 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_imm_packed = {_RANDOM_394[0], _RANDOM_393[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_csr_addr = _RANDOM_394[12:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_rob_idx = _RANDOM_394[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ldq_idx = _RANDOM_394[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stq_idx = _RANDOM_394[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_brob_idx = _RANDOM_394[31:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_395 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_pdst = _RANDOM_395[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_pop1 = _RANDOM_395[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_pop2 = _RANDOM_395[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_pop3 = _RANDOM_395[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_prs1_busy = _RANDOM_395[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_prs2_busy = _RANDOM_395[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_prs3_busy = _RANDOM_395[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_396 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_stale_pdst = {_RANDOM_396[5:0], _RANDOM_395[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_exception = _RANDOM_396[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_397 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_398 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_exc_cause = {_RANDOM_398[6:0], _RANDOM_397, _RANDOM_396[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_bypassable = _RANDOM_398[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_mem_cmd = _RANDOM_398[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_mem_typ = _RANDOM_398[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_fence = _RANDOM_398[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_fencei = _RANDOM_398[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_store = _RANDOM_398[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_amo = _RANDOM_398[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_load = _RANDOM_398[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_is_unique = _RANDOM_398[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_flush_on_commit = _RANDOM_398[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ldst = _RANDOM_398[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_399 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_lrs1 = {_RANDOM_399[1:0], _RANDOM_398[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_lrs2 = _RANDOM_399[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_lrs3 = _RANDOM_399[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_ldst_val = _RANDOM_399[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_dst_rtype = _RANDOM_399[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_lrs1_rtype = _RANDOM_399[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_lrs2_rtype = _RANDOM_399[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_frs3_en = _RANDOM_399[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_fp_val = _RANDOM_399[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_fp_single = _RANDOM_399[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_xcpt_if = _RANDOM_399[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_replay_if = _RANDOM_399[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_400 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_401 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_debug_wdata = {_RANDOM_401[25:0], _RANDOM_400, _RANDOM_399[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_402 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_10_debug_events_fetch_seq = {_RANDOM_402[25:0], _RANDOM_401[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_valid = _RANDOM_402[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_iw_state = _RANDOM_402[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_403 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_uopc = {_RANDOM_403[5:0], _RANDOM_402[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_404 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_inst = {_RANDOM_404[5:0], _RANDOM_403[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_405 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_pc = {_RANDOM_405[13:0], _RANDOM_404[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_fu_code = _RANDOM_405[21:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_br_type = _RANDOM_405[25:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_op1_sel = _RANDOM_405[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_op2_sel = _RANDOM_405[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_406 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_imm_sel = {_RANDOM_406[1:0], _RANDOM_405[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_op_fcn = _RANDOM_406[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_fcn_dw = _RANDOM_406[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_rf_wen = _RANDOM_406[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_csr_cmd = _RANDOM_406[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_is_load = _RANDOM_406[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_is_sta = _RANDOM_406[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ctrl_is_std = _RANDOM_406[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_wakeup_delay = _RANDOM_406[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_allocate_brtag = _RANDOM_406[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_br_or_jmp = _RANDOM_406[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_jump = _RANDOM_406[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_jal = _RANDOM_406[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_ret = _RANDOM_406[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_call = _RANDOM_406[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_mask = _RANDOM_406[29:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_407 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_tag = {_RANDOM_407[0], _RANDOM_406[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_prediction_bpd_predict_val = _RANDOM_407[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_prediction_bpd_predict_taken = _RANDOM_407[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_prediction_btb_hit = _RANDOM_407[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_prediction_btb_predicted = _RANDOM_407[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_br_prediction_is_br_or_jalr = _RANDOM_407[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stat_brjmp_mispredicted = _RANDOM_407[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stat_btb_made_pred = _RANDOM_407[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stat_btb_mispredicted = _RANDOM_407[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stat_bpd_made_pred = _RANDOM_407[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stat_bpd_mispredicted = _RANDOM_407[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_fetch_pc_lob = _RANDOM_407[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_408 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_imm_packed = {_RANDOM_408[1:0], _RANDOM_407[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_csr_addr = _RANDOM_408[13:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_rob_idx = _RANDOM_408[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ldq_idx = _RANDOM_408[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stq_idx = _RANDOM_408[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_409 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_brob_idx = {_RANDOM_409[0], _RANDOM_408[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_pdst = _RANDOM_409[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_pop1 = _RANDOM_409[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_pop2 = _RANDOM_409[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_pop3 = _RANDOM_409[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_prs1_busy = _RANDOM_409[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_prs2_busy = _RANDOM_409[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_prs3_busy = _RANDOM_409[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_410 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_stale_pdst = _RANDOM_410[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_exception = _RANDOM_410[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_411 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_412 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_exc_cause = {_RANDOM_412[7:0], _RANDOM_411, _RANDOM_410[31:8]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_bypassable = _RANDOM_412[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_mem_cmd = _RANDOM_412[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_mem_typ = _RANDOM_412[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_fence = _RANDOM_412[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_fencei = _RANDOM_412[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_store = _RANDOM_412[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_amo = _RANDOM_412[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_load = _RANDOM_412[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_is_unique = _RANDOM_412[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_flush_on_commit = _RANDOM_412[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ldst = _RANDOM_412[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_413 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_lrs1 = {_RANDOM_413[2:0], _RANDOM_412[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_lrs2 = _RANDOM_413[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_lrs3 = _RANDOM_413[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_ldst_val = _RANDOM_413[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_dst_rtype = _RANDOM_413[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_lrs1_rtype = _RANDOM_413[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_lrs2_rtype = _RANDOM_413[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_frs3_en = _RANDOM_413[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_fp_val = _RANDOM_413[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_fp_single = _RANDOM_413[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_xcpt_if = _RANDOM_413[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_replay_if = _RANDOM_413[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_414 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_415 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_debug_wdata = {_RANDOM_415[26:0], _RANDOM_414, _RANDOM_413[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_416 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_11_debug_events_fetch_seq = {_RANDOM_416[26:0], _RANDOM_415[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_valid = _RANDOM_416[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_iw_state = _RANDOM_416[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_417 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_uopc = {_RANDOM_417[6:0], _RANDOM_416[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_418 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_inst = {_RANDOM_418[6:0], _RANDOM_417[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_419 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_pc = {_RANDOM_419[14:0], _RANDOM_418[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_fu_code = _RANDOM_419[22:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_br_type = _RANDOM_419[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_op1_sel = _RANDOM_419[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_op2_sel = _RANDOM_419[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_420 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_imm_sel = _RANDOM_420[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_op_fcn = _RANDOM_420[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_fcn_dw = _RANDOM_420[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_rf_wen = _RANDOM_420[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_csr_cmd = _RANDOM_420[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_is_load = _RANDOM_420[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_is_sta = _RANDOM_420[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ctrl_is_std = _RANDOM_420[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_wakeup_delay = _RANDOM_420[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_allocate_brtag = _RANDOM_420[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_br_or_jmp = _RANDOM_420[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_jump = _RANDOM_420[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_jal = _RANDOM_420[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_ret = _RANDOM_420[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_call = _RANDOM_420[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_mask = _RANDOM_420[30:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_421 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_tag = {_RANDOM_421[1:0], _RANDOM_420[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_prediction_bpd_predict_val = _RANDOM_421[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_prediction_bpd_predict_taken = _RANDOM_421[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_prediction_btb_hit = _RANDOM_421[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_prediction_btb_predicted = _RANDOM_421[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_br_prediction_is_br_or_jalr = _RANDOM_421[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stat_brjmp_mispredicted = _RANDOM_421[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stat_btb_made_pred = _RANDOM_421[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stat_btb_mispredicted = _RANDOM_421[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stat_bpd_made_pred = _RANDOM_421[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stat_bpd_mispredicted = _RANDOM_421[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_fetch_pc_lob = _RANDOM_421[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_422 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_imm_packed = {_RANDOM_422[2:0], _RANDOM_421[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_csr_addr = _RANDOM_422[14:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_rob_idx = _RANDOM_422[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ldq_idx = _RANDOM_422[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stq_idx = _RANDOM_422[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_423 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_brob_idx = {_RANDOM_423[1:0], _RANDOM_422[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_pdst = _RANDOM_423[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_pop1 = _RANDOM_423[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_pop2 = _RANDOM_423[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_pop3 = _RANDOM_423[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_prs1_busy = _RANDOM_423[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_prs2_busy = _RANDOM_423[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_424 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_prs3_busy = _RANDOM_424[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_stale_pdst = _RANDOM_424[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_exception = _RANDOM_424[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_425 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_426 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_exc_cause = {_RANDOM_426[8:0], _RANDOM_425, _RANDOM_424[31:9]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_bypassable = _RANDOM_426[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_mem_cmd = _RANDOM_426[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_mem_typ = _RANDOM_426[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_fence = _RANDOM_426[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_fencei = _RANDOM_426[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_store = _RANDOM_426[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_amo = _RANDOM_426[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_load = _RANDOM_426[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_is_unique = _RANDOM_426[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_flush_on_commit = _RANDOM_426[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ldst = _RANDOM_426[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_427 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_lrs1 = {_RANDOM_427[3:0], _RANDOM_426[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_lrs2 = _RANDOM_427[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_lrs3 = _RANDOM_427[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_ldst_val = _RANDOM_427[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_dst_rtype = _RANDOM_427[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_lrs1_rtype = _RANDOM_427[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_lrs2_rtype = _RANDOM_427[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_frs3_en = _RANDOM_427[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_fp_val = _RANDOM_427[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_fp_single = _RANDOM_427[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_xcpt_if = _RANDOM_427[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_replay_if = _RANDOM_427[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_428 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_429 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_debug_wdata = {_RANDOM_429[27:0], _RANDOM_428, _RANDOM_427[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_430 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_12_debug_events_fetch_seq = {_RANDOM_430[27:0], _RANDOM_429[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_valid = _RANDOM_430[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_iw_state = _RANDOM_430[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_431 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_uopc = {_RANDOM_431[7:0], _RANDOM_430[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_432 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_inst = {_RANDOM_432[7:0], _RANDOM_431[31:8]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_433 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_pc = {_RANDOM_433[15:0], _RANDOM_432[31:8]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_fu_code = _RANDOM_433[23:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_br_type = _RANDOM_433[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_op1_sel = _RANDOM_433[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_434 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_op2_sel = {_RANDOM_434[0], _RANDOM_433[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_imm_sel = _RANDOM_434[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_op_fcn = _RANDOM_434[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_fcn_dw = _RANDOM_434[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_rf_wen = _RANDOM_434[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_csr_cmd = _RANDOM_434[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_is_load = _RANDOM_434[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_is_sta = _RANDOM_434[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ctrl_is_std = _RANDOM_434[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_wakeup_delay = _RANDOM_434[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_allocate_brtag = _RANDOM_434[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_br_or_jmp = _RANDOM_434[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_jump = _RANDOM_434[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_jal = _RANDOM_434[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_ret = _RANDOM_434[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_call = _RANDOM_434[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_mask = _RANDOM_434[31:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_435 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_tag = _RANDOM_435[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_prediction_bpd_predict_val = _RANDOM_435[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_prediction_bpd_predict_taken = _RANDOM_435[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_prediction_btb_hit = _RANDOM_435[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_prediction_btb_predicted = _RANDOM_435[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_br_prediction_is_br_or_jalr = _RANDOM_435[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stat_brjmp_mispredicted = _RANDOM_435[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stat_btb_made_pred = _RANDOM_435[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stat_btb_mispredicted = _RANDOM_435[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stat_bpd_made_pred = _RANDOM_435[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stat_bpd_mispredicted = _RANDOM_435[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_fetch_pc_lob = _RANDOM_435[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_436 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_imm_packed = {_RANDOM_436[3:0], _RANDOM_435[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_csr_addr = _RANDOM_436[15:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_rob_idx = _RANDOM_436[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ldq_idx = _RANDOM_436[25:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stq_idx = _RANDOM_436[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_437 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_brob_idx = {_RANDOM_437[2:0], _RANDOM_436[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_pdst = _RANDOM_437[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_pop1 = _RANDOM_437[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_pop2 = _RANDOM_437[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_pop3 = _RANDOM_437[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_prs1_busy = _RANDOM_437[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_438 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_prs2_busy = _RANDOM_438[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_prs3_busy = _RANDOM_438[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_stale_pdst = _RANDOM_438[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_exception = _RANDOM_438[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_439 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_440 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_exc_cause = {_RANDOM_440[9:0], _RANDOM_439, _RANDOM_438[31:10]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_bypassable = _RANDOM_440[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_mem_cmd = _RANDOM_440[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_mem_typ = _RANDOM_440[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_fence = _RANDOM_440[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_fencei = _RANDOM_440[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_store = _RANDOM_440[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_amo = _RANDOM_440[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_load = _RANDOM_440[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_is_unique = _RANDOM_440[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_flush_on_commit = _RANDOM_440[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ldst = _RANDOM_440[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_441 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_lrs1 = {_RANDOM_441[4:0], _RANDOM_440[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_lrs2 = _RANDOM_441[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_lrs3 = _RANDOM_441[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_ldst_val = _RANDOM_441[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_dst_rtype = _RANDOM_441[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_lrs1_rtype = _RANDOM_441[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_lrs2_rtype = _RANDOM_441[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_frs3_en = _RANDOM_441[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_fp_val = _RANDOM_441[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_fp_single = _RANDOM_441[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_xcpt_if = _RANDOM_441[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_replay_if = _RANDOM_441[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_442 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_443 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_debug_wdata = {_RANDOM_443[28:0], _RANDOM_442, _RANDOM_441[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_444 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_13_debug_events_fetch_seq = {_RANDOM_444[28:0], _RANDOM_443[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_valid = _RANDOM_444[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_iw_state = _RANDOM_444[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_445 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_uopc = _RANDOM_445[8:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_446 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_inst = {_RANDOM_446[8:0], _RANDOM_445[31:9]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_447 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_pc = {_RANDOM_447[16:0], _RANDOM_446[31:9]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_fu_code = _RANDOM_447[24:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_br_type = _RANDOM_447[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_op1_sel = _RANDOM_447[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_448 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_op2_sel = {_RANDOM_448[1:0], _RANDOM_447[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_imm_sel = _RANDOM_448[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_op_fcn = _RANDOM_448[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_fcn_dw = _RANDOM_448[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_rf_wen = _RANDOM_448[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_csr_cmd = _RANDOM_448[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_is_load = _RANDOM_448[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_is_sta = _RANDOM_448[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ctrl_is_std = _RANDOM_448[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_wakeup_delay = _RANDOM_448[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_allocate_brtag = _RANDOM_448[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_br_or_jmp = _RANDOM_448[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_jump = _RANDOM_448[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_jal = _RANDOM_448[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_ret = _RANDOM_448[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_call = _RANDOM_448[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_449 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_mask = {_RANDOM_449[0], _RANDOM_448[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_tag = _RANDOM_449[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_prediction_bpd_predict_val = _RANDOM_449[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_prediction_bpd_predict_taken = _RANDOM_449[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_prediction_btb_hit = _RANDOM_449[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_prediction_btb_predicted = _RANDOM_449[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_br_prediction_is_br_or_jalr = _RANDOM_449[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stat_brjmp_mispredicted = _RANDOM_449[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stat_btb_made_pred = _RANDOM_449[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stat_btb_mispredicted = _RANDOM_449[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stat_bpd_made_pred = _RANDOM_449[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stat_bpd_mispredicted = _RANDOM_449[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_fetch_pc_lob = _RANDOM_449[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_450 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_imm_packed = {_RANDOM_450[4:0], _RANDOM_449[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_csr_addr = _RANDOM_450[16:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_rob_idx = _RANDOM_450[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ldq_idx = _RANDOM_450[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stq_idx = _RANDOM_450[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_451 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_brob_idx = {_RANDOM_451[3:0], _RANDOM_450[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_pdst = _RANDOM_451[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_pop1 = _RANDOM_451[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_pop2 = _RANDOM_451[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_pop3 = _RANDOM_451[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_452 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_prs1_busy = _RANDOM_452[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_prs2_busy = _RANDOM_452[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_prs3_busy = _RANDOM_452[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_stale_pdst = _RANDOM_452[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_exception = _RANDOM_452[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_453 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_454 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_exc_cause = {_RANDOM_454[10:0], _RANDOM_453, _RANDOM_452[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_bypassable = _RANDOM_454[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_mem_cmd = _RANDOM_454[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_mem_typ = _RANDOM_454[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_fence = _RANDOM_454[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_fencei = _RANDOM_454[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_store = _RANDOM_454[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_amo = _RANDOM_454[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_load = _RANDOM_454[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_is_unique = _RANDOM_454[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_flush_on_commit = _RANDOM_454[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ldst = _RANDOM_454[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_455 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_lrs1 = _RANDOM_455[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_lrs2 = _RANDOM_455[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_lrs3 = _RANDOM_455[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_ldst_val = _RANDOM_455[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_dst_rtype = _RANDOM_455[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_lrs1_rtype = _RANDOM_455[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_lrs2_rtype = _RANDOM_455[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_frs3_en = _RANDOM_455[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_fp_val = _RANDOM_455[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_fp_single = _RANDOM_455[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_xcpt_if = _RANDOM_455[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_replay_if = _RANDOM_455[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_456 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_457 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_debug_wdata = {_RANDOM_457[29:0], _RANDOM_456, _RANDOM_455[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_458 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_14_debug_events_fetch_seq = {_RANDOM_458[29:0], _RANDOM_457[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_valid = _RANDOM_458[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_459 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_iw_state = {_RANDOM_459[0], _RANDOM_458[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_uopc = _RANDOM_459[9:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_460 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_inst = {_RANDOM_460[9:0], _RANDOM_459[31:10]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_461 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_pc = {_RANDOM_461[17:0], _RANDOM_460[31:10]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_fu_code = _RANDOM_461[25:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_br_type = _RANDOM_461[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_op1_sel = _RANDOM_461[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_462 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_op2_sel = _RANDOM_462[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_imm_sel = _RANDOM_462[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_op_fcn = _RANDOM_462[9:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_fcn_dw = _RANDOM_462[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_rf_wen = _RANDOM_462[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_csr_cmd = _RANDOM_462[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_is_load = _RANDOM_462[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_is_sta = _RANDOM_462[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ctrl_is_std = _RANDOM_462[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_wakeup_delay = _RANDOM_462[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_allocate_brtag = _RANDOM_462[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_br_or_jmp = _RANDOM_462[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_jump = _RANDOM_462[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_jal = _RANDOM_462[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_ret = _RANDOM_462[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_call = _RANDOM_462[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_463 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_mask = {_RANDOM_463[1:0], _RANDOM_462[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_tag = _RANDOM_463[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_prediction_bpd_predict_val = _RANDOM_463[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_prediction_bpd_predict_taken = _RANDOM_463[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_prediction_btb_hit = _RANDOM_463[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_prediction_btb_predicted = _RANDOM_463[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_br_prediction_is_br_or_jalr = _RANDOM_463[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stat_brjmp_mispredicted = _RANDOM_463[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stat_btb_made_pred = _RANDOM_463[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stat_btb_mispredicted = _RANDOM_463[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stat_bpd_made_pred = _RANDOM_463[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stat_bpd_mispredicted = _RANDOM_463[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_fetch_pc_lob = _RANDOM_463[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_464 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_imm_packed = {_RANDOM_464[5:0], _RANDOM_463[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_csr_addr = _RANDOM_464[17:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_rob_idx = _RANDOM_464[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ldq_idx = _RANDOM_464[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stq_idx = _RANDOM_464[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_465 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_brob_idx = _RANDOM_465[4:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_pdst = _RANDOM_465[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_pop1 = _RANDOM_465[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_pop2 = _RANDOM_465[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_466 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_pop3 = {_RANDOM_466[0], _RANDOM_465[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_prs1_busy = _RANDOM_466[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_prs2_busy = _RANDOM_466[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_prs3_busy = _RANDOM_466[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_stale_pdst = _RANDOM_466[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_exception = _RANDOM_466[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_467 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_468 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_exc_cause = {_RANDOM_468[11:0], _RANDOM_467, _RANDOM_466[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_bypassable = _RANDOM_468[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_mem_cmd = _RANDOM_468[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_mem_typ = _RANDOM_468[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_fence = _RANDOM_468[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_fencei = _RANDOM_468[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_store = _RANDOM_468[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_amo = _RANDOM_468[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_load = _RANDOM_468[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_is_unique = _RANDOM_468[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_flush_on_commit = _RANDOM_468[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_469 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ldst = {_RANDOM_469[0], _RANDOM_468[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_lrs1 = _RANDOM_469[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_lrs2 = _RANDOM_469[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_lrs3 = _RANDOM_469[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_ldst_val = _RANDOM_469[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_dst_rtype = _RANDOM_469[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_lrs1_rtype = _RANDOM_469[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_lrs2_rtype = _RANDOM_469[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_frs3_en = _RANDOM_469[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_fp_val = _RANDOM_469[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_fp_single = _RANDOM_469[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_xcpt_if = _RANDOM_469[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_replay_if = _RANDOM_469[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_470 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_471 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_debug_wdata = {_RANDOM_471[30:0], _RANDOM_470, _RANDOM_469[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_472 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_15_debug_events_fetch_seq = {_RANDOM_472[30:0], _RANDOM_471[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_valid = _RANDOM_472[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_473 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_iw_state = _RANDOM_473[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_uopc = _RANDOM_473[10:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_474 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_inst = {_RANDOM_474[10:0], _RANDOM_473[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_475 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_pc = {_RANDOM_475[18:0], _RANDOM_474[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_fu_code = _RANDOM_475[26:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_br_type = _RANDOM_475[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_476 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_op1_sel = {_RANDOM_476[0], _RANDOM_475[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_op2_sel = _RANDOM_476[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_imm_sel = _RANDOM_476[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_op_fcn = _RANDOM_476[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_fcn_dw = _RANDOM_476[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_rf_wen = _RANDOM_476[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_csr_cmd = _RANDOM_476[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_is_load = _RANDOM_476[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_is_sta = _RANDOM_476[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ctrl_is_std = _RANDOM_476[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_wakeup_delay = _RANDOM_476[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_allocate_brtag = _RANDOM_476[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_br_or_jmp = _RANDOM_476[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_jump = _RANDOM_476[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_jal = _RANDOM_476[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_ret = _RANDOM_476[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_call = _RANDOM_476[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_477 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_mask = {_RANDOM_477[2:0], _RANDOM_476[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_tag = _RANDOM_477[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_prediction_bpd_predict_val = _RANDOM_477[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_prediction_bpd_predict_taken = _RANDOM_477[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_prediction_btb_hit = _RANDOM_477[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_prediction_btb_predicted = _RANDOM_477[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_br_prediction_is_br_or_jalr = _RANDOM_477[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stat_brjmp_mispredicted = _RANDOM_477[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stat_btb_made_pred = _RANDOM_477[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stat_btb_mispredicted = _RANDOM_477[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stat_bpd_made_pred = _RANDOM_477[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stat_bpd_mispredicted = _RANDOM_477[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_fetch_pc_lob = _RANDOM_477[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_478 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_imm_packed = {_RANDOM_478[6:0], _RANDOM_477[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_csr_addr = _RANDOM_478[18:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_rob_idx = _RANDOM_478[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ldq_idx = _RANDOM_478[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_479 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stq_idx = {_RANDOM_479[0], _RANDOM_478[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_brob_idx = _RANDOM_479[5:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_pdst = _RANDOM_479[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_pop1 = _RANDOM_479[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_pop2 = _RANDOM_479[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_480 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_pop3 = {_RANDOM_480[1:0], _RANDOM_479[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_prs1_busy = _RANDOM_480[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_prs2_busy = _RANDOM_480[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_prs3_busy = _RANDOM_480[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_stale_pdst = _RANDOM_480[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_exception = _RANDOM_480[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_481 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_482 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_exc_cause = {_RANDOM_482[12:0], _RANDOM_481, _RANDOM_480[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_bypassable = _RANDOM_482[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_mem_cmd = _RANDOM_482[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_mem_typ = _RANDOM_482[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_fence = _RANDOM_482[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_fencei = _RANDOM_482[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_store = _RANDOM_482[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_amo = _RANDOM_482[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_load = _RANDOM_482[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_is_unique = _RANDOM_482[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_flush_on_commit = _RANDOM_482[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_483 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ldst = {_RANDOM_483[1:0], _RANDOM_482[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_lrs1 = _RANDOM_483[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_lrs2 = _RANDOM_483[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_lrs3 = _RANDOM_483[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_ldst_val = _RANDOM_483[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_dst_rtype = _RANDOM_483[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_lrs1_rtype = _RANDOM_483[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_lrs2_rtype = _RANDOM_483[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_frs3_en = _RANDOM_483[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_fp_val = _RANDOM_483[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_fp_single = _RANDOM_483[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_xcpt_if = _RANDOM_483[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_replay_if = _RANDOM_483[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_484 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_485 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_debug_wdata = {_RANDOM_485, _RANDOM_484};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_486 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_16_debug_events_fetch_seq = _RANDOM_486;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_487 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_valid = _RANDOM_487[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_iw_state = _RANDOM_487[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_uopc = _RANDOM_487[11:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_488 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_inst = {_RANDOM_488[11:0], _RANDOM_487[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_489 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_pc = {_RANDOM_489[19:0], _RANDOM_488[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_fu_code = _RANDOM_489[27:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_br_type = _RANDOM_489[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_490 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_op1_sel = _RANDOM_490[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_op2_sel = _RANDOM_490[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_imm_sel = _RANDOM_490[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_op_fcn = _RANDOM_490[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_fcn_dw = _RANDOM_490[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_rf_wen = _RANDOM_490[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_csr_cmd = _RANDOM_490[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_is_load = _RANDOM_490[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_is_sta = _RANDOM_490[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ctrl_is_std = _RANDOM_490[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_wakeup_delay = _RANDOM_490[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_allocate_brtag = _RANDOM_490[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_br_or_jmp = _RANDOM_490[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_jump = _RANDOM_490[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_jal = _RANDOM_490[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_ret = _RANDOM_490[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_call = _RANDOM_490[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_491 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_mask = {_RANDOM_491[3:0], _RANDOM_490[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_tag = _RANDOM_491[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_prediction_bpd_predict_val = _RANDOM_491[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_prediction_bpd_predict_taken = _RANDOM_491[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_prediction_btb_hit = _RANDOM_491[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_prediction_btb_predicted = _RANDOM_491[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_br_prediction_is_br_or_jalr = _RANDOM_491[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stat_brjmp_mispredicted = _RANDOM_491[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stat_btb_made_pred = _RANDOM_491[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stat_btb_mispredicted = _RANDOM_491[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stat_bpd_made_pred = _RANDOM_491[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stat_bpd_mispredicted = _RANDOM_491[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_fetch_pc_lob = _RANDOM_491[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_492 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_imm_packed = {_RANDOM_492[7:0], _RANDOM_491[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_csr_addr = _RANDOM_492[19:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_rob_idx = _RANDOM_492[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ldq_idx = _RANDOM_492[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_493 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stq_idx = {_RANDOM_493[1:0], _RANDOM_492[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_brob_idx = _RANDOM_493[6:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_pdst = _RANDOM_493[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_pop1 = _RANDOM_493[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_pop2 = _RANDOM_493[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_494 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_pop3 = {_RANDOM_494[2:0], _RANDOM_493[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_prs1_busy = _RANDOM_494[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_prs2_busy = _RANDOM_494[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_prs3_busy = _RANDOM_494[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_stale_pdst = _RANDOM_494[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_exception = _RANDOM_494[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_495 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_496 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_exc_cause = {_RANDOM_496[13:0], _RANDOM_495, _RANDOM_494[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_bypassable = _RANDOM_496[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_mem_cmd = _RANDOM_496[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_mem_typ = _RANDOM_496[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_fence = _RANDOM_496[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_fencei = _RANDOM_496[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_store = _RANDOM_496[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_amo = _RANDOM_496[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_load = _RANDOM_496[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_is_unique = _RANDOM_496[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_flush_on_commit = _RANDOM_496[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_497 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ldst = {_RANDOM_497[2:0], _RANDOM_496[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_lrs1 = _RANDOM_497[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_lrs2 = _RANDOM_497[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_lrs3 = _RANDOM_497[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_ldst_val = _RANDOM_497[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_dst_rtype = _RANDOM_497[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_lrs1_rtype = _RANDOM_497[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_lrs2_rtype = _RANDOM_497[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_frs3_en = _RANDOM_497[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_fp_val = _RANDOM_497[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_fp_single = _RANDOM_497[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_xcpt_if = _RANDOM_497[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_498 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_replay_if = _RANDOM_498[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_499 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_500 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_debug_wdata = {_RANDOM_500[0], _RANDOM_499, _RANDOM_498[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_501 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_17_debug_events_fetch_seq = {_RANDOM_501[0], _RANDOM_500[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_valid = _RANDOM_501[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_iw_state = _RANDOM_501[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_uopc = _RANDOM_501[12:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_502 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_inst = {_RANDOM_502[12:0], _RANDOM_501[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_503 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_pc = {_RANDOM_503[20:0], _RANDOM_502[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_fu_code = _RANDOM_503[28:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_504 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_br_type = {_RANDOM_504[0], _RANDOM_503[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_op1_sel = _RANDOM_504[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_op2_sel = _RANDOM_504[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_imm_sel = _RANDOM_504[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_op_fcn = _RANDOM_504[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_fcn_dw = _RANDOM_504[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_rf_wen = _RANDOM_504[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_csr_cmd = _RANDOM_504[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_is_load = _RANDOM_504[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_is_sta = _RANDOM_504[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ctrl_is_std = _RANDOM_504[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_wakeup_delay = _RANDOM_504[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_allocate_brtag = _RANDOM_504[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_br_or_jmp = _RANDOM_504[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_jump = _RANDOM_504[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_jal = _RANDOM_504[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_ret = _RANDOM_504[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_call = _RANDOM_504[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_505 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_mask = {_RANDOM_505[4:0], _RANDOM_504[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_tag = _RANDOM_505[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_prediction_bpd_predict_val = _RANDOM_505[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_prediction_bpd_predict_taken = _RANDOM_505[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_prediction_btb_hit = _RANDOM_505[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_prediction_btb_predicted = _RANDOM_505[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_br_prediction_is_br_or_jalr = _RANDOM_505[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stat_brjmp_mispredicted = _RANDOM_505[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stat_btb_made_pred = _RANDOM_505[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stat_btb_mispredicted = _RANDOM_505[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stat_bpd_made_pred = _RANDOM_505[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stat_bpd_mispredicted = _RANDOM_505[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_fetch_pc_lob = _RANDOM_505[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_506 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_imm_packed = {_RANDOM_506[8:0], _RANDOM_505[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_csr_addr = _RANDOM_506[20:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_rob_idx = _RANDOM_506[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ldq_idx = _RANDOM_506[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_507 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stq_idx = {_RANDOM_507[2:0], _RANDOM_506[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_brob_idx = _RANDOM_507[7:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_pdst = _RANDOM_507[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_pop1 = _RANDOM_507[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_pop2 = _RANDOM_507[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_508 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_pop3 = {_RANDOM_508[3:0], _RANDOM_507[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_prs1_busy = _RANDOM_508[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_prs2_busy = _RANDOM_508[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_prs3_busy = _RANDOM_508[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_stale_pdst = _RANDOM_508[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_exception = _RANDOM_508[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_509 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_510 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_exc_cause = {_RANDOM_510[14:0], _RANDOM_509, _RANDOM_508[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_bypassable = _RANDOM_510[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_mem_cmd = _RANDOM_510[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_mem_typ = _RANDOM_510[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_fence = _RANDOM_510[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_fencei = _RANDOM_510[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_store = _RANDOM_510[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_amo = _RANDOM_510[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_load = _RANDOM_510[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_is_unique = _RANDOM_510[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_flush_on_commit = _RANDOM_510[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_511 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ldst = {_RANDOM_511[3:0], _RANDOM_510[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_lrs1 = _RANDOM_511[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_lrs2 = _RANDOM_511[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_lrs3 = _RANDOM_511[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_ldst_val = _RANDOM_511[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_dst_rtype = _RANDOM_511[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_lrs1_rtype = _RANDOM_511[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_lrs2_rtype = _RANDOM_511[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_frs3_en = _RANDOM_511[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_fp_val = _RANDOM_511[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_fp_single = _RANDOM_511[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_512 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_xcpt_if = _RANDOM_512[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_replay_if = _RANDOM_512[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_513 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_514 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_debug_wdata = {_RANDOM_514[1:0], _RANDOM_513, _RANDOM_512[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_515 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_18_debug_events_fetch_seq = {_RANDOM_515[1:0], _RANDOM_514[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_valid = _RANDOM_515[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_iw_state = _RANDOM_515[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_uopc = _RANDOM_515[13:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_516 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_inst = {_RANDOM_516[13:0], _RANDOM_515[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_517 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_pc = {_RANDOM_517[21:0], _RANDOM_516[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_fu_code = _RANDOM_517[29:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_518 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_br_type = {_RANDOM_518[1:0], _RANDOM_517[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_op1_sel = _RANDOM_518[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_op2_sel = _RANDOM_518[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_imm_sel = _RANDOM_518[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_op_fcn = _RANDOM_518[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_fcn_dw = _RANDOM_518[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_rf_wen = _RANDOM_518[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_csr_cmd = _RANDOM_518[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_is_load = _RANDOM_518[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_is_sta = _RANDOM_518[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ctrl_is_std = _RANDOM_518[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_wakeup_delay = _RANDOM_518[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_allocate_brtag = _RANDOM_518[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_br_or_jmp = _RANDOM_518[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_jump = _RANDOM_518[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_jal = _RANDOM_518[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_ret = _RANDOM_518[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_call = _RANDOM_518[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_519 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_mask = {_RANDOM_519[5:0], _RANDOM_518[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_tag = _RANDOM_519[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_prediction_bpd_predict_val = _RANDOM_519[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_prediction_bpd_predict_taken = _RANDOM_519[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_prediction_btb_hit = _RANDOM_519[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_prediction_btb_predicted = _RANDOM_519[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_br_prediction_is_br_or_jalr = _RANDOM_519[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stat_brjmp_mispredicted = _RANDOM_519[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stat_btb_made_pred = _RANDOM_519[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stat_btb_mispredicted = _RANDOM_519[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stat_bpd_made_pred = _RANDOM_519[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stat_bpd_mispredicted = _RANDOM_519[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_fetch_pc_lob = _RANDOM_519[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_520 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_imm_packed = {_RANDOM_520[9:0], _RANDOM_519[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_csr_addr = _RANDOM_520[21:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_rob_idx = _RANDOM_520[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ldq_idx = _RANDOM_520[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_521 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stq_idx = _RANDOM_521[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_brob_idx = _RANDOM_521[8:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_pdst = _RANDOM_521[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_pop1 = _RANDOM_521[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_pop2 = _RANDOM_521[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_522 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_pop3 = {_RANDOM_522[4:0], _RANDOM_521[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_prs1_busy = _RANDOM_522[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_prs2_busy = _RANDOM_522[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_prs3_busy = _RANDOM_522[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_stale_pdst = _RANDOM_522[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_exception = _RANDOM_522[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_523 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_524 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_exc_cause = {_RANDOM_524[15:0], _RANDOM_523, _RANDOM_522[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_bypassable = _RANDOM_524[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_mem_cmd = _RANDOM_524[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_mem_typ = _RANDOM_524[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_fence = _RANDOM_524[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_fencei = _RANDOM_524[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_store = _RANDOM_524[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_amo = _RANDOM_524[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_load = _RANDOM_524[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_is_unique = _RANDOM_524[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_flush_on_commit = _RANDOM_524[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_525 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ldst = {_RANDOM_525[4:0], _RANDOM_524[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_lrs1 = _RANDOM_525[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_lrs2 = _RANDOM_525[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_lrs3 = _RANDOM_525[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_ldst_val = _RANDOM_525[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_dst_rtype = _RANDOM_525[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_lrs1_rtype = _RANDOM_525[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_lrs2_rtype = _RANDOM_525[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_frs3_en = _RANDOM_525[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_fp_val = _RANDOM_525[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_526 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_fp_single = _RANDOM_526[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_xcpt_if = _RANDOM_526[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_replay_if = _RANDOM_526[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_527 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_528 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_debug_wdata = {_RANDOM_528[2:0], _RANDOM_527, _RANDOM_526[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_529 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_19_debug_events_fetch_seq = {_RANDOM_529[2:0], _RANDOM_528[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_valid = _RANDOM_529[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_iw_state = _RANDOM_529[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_uopc = _RANDOM_529[14:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_530 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_inst = {_RANDOM_530[14:0], _RANDOM_529[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_531 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_pc = {_RANDOM_531[22:0], _RANDOM_530[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_fu_code = _RANDOM_531[30:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_532 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_br_type = {_RANDOM_532[2:0], _RANDOM_531[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_op1_sel = _RANDOM_532[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_op2_sel = _RANDOM_532[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_imm_sel = _RANDOM_532[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_op_fcn = _RANDOM_532[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_fcn_dw = _RANDOM_532[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_rf_wen = _RANDOM_532[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_csr_cmd = _RANDOM_532[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_is_load = _RANDOM_532[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_is_sta = _RANDOM_532[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ctrl_is_std = _RANDOM_532[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_wakeup_delay = _RANDOM_532[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_allocate_brtag = _RANDOM_532[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_br_or_jmp = _RANDOM_532[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_jump = _RANDOM_532[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_jal = _RANDOM_532[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_ret = _RANDOM_532[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_call = _RANDOM_532[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_533 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_mask = {_RANDOM_533[6:0], _RANDOM_532[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_tag = _RANDOM_533[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_prediction_bpd_predict_val = _RANDOM_533[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_prediction_bpd_predict_taken = _RANDOM_533[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_prediction_btb_hit = _RANDOM_533[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_prediction_btb_predicted = _RANDOM_533[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_br_prediction_is_br_or_jalr = _RANDOM_533[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stat_brjmp_mispredicted = _RANDOM_533[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stat_btb_made_pred = _RANDOM_533[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stat_btb_mispredicted = _RANDOM_533[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stat_bpd_made_pred = _RANDOM_533[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stat_bpd_mispredicted = _RANDOM_533[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_fetch_pc_lob = _RANDOM_533[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_534 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_imm_packed = {_RANDOM_534[10:0], _RANDOM_533[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_csr_addr = _RANDOM_534[22:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_rob_idx = _RANDOM_534[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_535 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ldq_idx = {_RANDOM_535[0], _RANDOM_534[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stq_idx = _RANDOM_535[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_brob_idx = _RANDOM_535[9:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_pdst = _RANDOM_535[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_pop1 = _RANDOM_535[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_pop2 = _RANDOM_535[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_536 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_pop3 = {_RANDOM_536[5:0], _RANDOM_535[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_prs1_busy = _RANDOM_536[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_prs2_busy = _RANDOM_536[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_prs3_busy = _RANDOM_536[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_stale_pdst = _RANDOM_536[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_exception = _RANDOM_536[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_537 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_538 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_exc_cause = {_RANDOM_538[16:0], _RANDOM_537, _RANDOM_536[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_bypassable = _RANDOM_538[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_mem_cmd = _RANDOM_538[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_mem_typ = _RANDOM_538[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_fence = _RANDOM_538[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_fencei = _RANDOM_538[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_store = _RANDOM_538[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_amo = _RANDOM_538[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_load = _RANDOM_538[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_is_unique = _RANDOM_538[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_flush_on_commit = _RANDOM_538[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_539 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ldst = _RANDOM_539[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_lrs1 = _RANDOM_539[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_lrs2 = _RANDOM_539[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_lrs3 = _RANDOM_539[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_ldst_val = _RANDOM_539[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_dst_rtype = _RANDOM_539[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_lrs1_rtype = _RANDOM_539[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_lrs2_rtype = _RANDOM_539[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_frs3_en = _RANDOM_539[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_540 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_fp_val = _RANDOM_540[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_fp_single = _RANDOM_540[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_xcpt_if = _RANDOM_540[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_replay_if = _RANDOM_540[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_541 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_542 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_debug_wdata = {_RANDOM_542[3:0], _RANDOM_541, _RANDOM_540[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_543 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_20_debug_events_fetch_seq = {_RANDOM_543[3:0], _RANDOM_542[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_valid = _RANDOM_543[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_iw_state = _RANDOM_543[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_uopc = _RANDOM_543[15:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_544 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_inst = {_RANDOM_544[15:0], _RANDOM_543[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_545 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_pc = {_RANDOM_545[23:0], _RANDOM_544[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_fu_code = _RANDOM_545[31:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_546 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_br_type = _RANDOM_546[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_op1_sel = _RANDOM_546[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_op2_sel = _RANDOM_546[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_imm_sel = _RANDOM_546[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_op_fcn = _RANDOM_546[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_fcn_dw = _RANDOM_546[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_rf_wen = _RANDOM_546[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_csr_cmd = _RANDOM_546[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_is_load = _RANDOM_546[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_is_sta = _RANDOM_546[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ctrl_is_std = _RANDOM_546[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_wakeup_delay = _RANDOM_546[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_allocate_brtag = _RANDOM_546[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_br_or_jmp = _RANDOM_546[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_jump = _RANDOM_546[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_jal = _RANDOM_546[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_ret = _RANDOM_546[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_call = _RANDOM_546[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_547 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_mask = _RANDOM_547[7:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_tag = _RANDOM_547[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_prediction_bpd_predict_val = _RANDOM_547[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_prediction_bpd_predict_taken = _RANDOM_547[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_prediction_btb_hit = _RANDOM_547[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_prediction_btb_predicted = _RANDOM_547[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_br_prediction_is_br_or_jalr = _RANDOM_547[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stat_brjmp_mispredicted = _RANDOM_547[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stat_btb_made_pred = _RANDOM_547[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stat_btb_mispredicted = _RANDOM_547[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stat_bpd_made_pred = _RANDOM_547[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stat_bpd_mispredicted = _RANDOM_547[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_fetch_pc_lob = _RANDOM_547[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_548 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_imm_packed = {_RANDOM_548[11:0], _RANDOM_547[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_csr_addr = _RANDOM_548[23:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_rob_idx = _RANDOM_548[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_549 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ldq_idx = {_RANDOM_549[1:0], _RANDOM_548[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stq_idx = _RANDOM_549[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_brob_idx = _RANDOM_549[10:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_pdst = _RANDOM_549[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_pop1 = _RANDOM_549[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_pop2 = _RANDOM_549[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_550 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_pop3 = _RANDOM_550[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_prs1_busy = _RANDOM_550[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_prs2_busy = _RANDOM_550[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_prs3_busy = _RANDOM_550[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_stale_pdst = _RANDOM_550[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_exception = _RANDOM_550[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_551 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_552 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_exc_cause = {_RANDOM_552[17:0], _RANDOM_551, _RANDOM_550[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_bypassable = _RANDOM_552[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_mem_cmd = _RANDOM_552[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_mem_typ = _RANDOM_552[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_fence = _RANDOM_552[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_fencei = _RANDOM_552[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_store = _RANDOM_552[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_amo = _RANDOM_552[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_load = _RANDOM_552[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_is_unique = _RANDOM_552[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_553 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_flush_on_commit = _RANDOM_553[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ldst = _RANDOM_553[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_lrs1 = _RANDOM_553[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_lrs2 = _RANDOM_553[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_lrs3 = _RANDOM_553[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_ldst_val = _RANDOM_553[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_dst_rtype = _RANDOM_553[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_lrs1_rtype = _RANDOM_553[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_lrs2_rtype = _RANDOM_553[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_554 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_frs3_en = _RANDOM_554[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_fp_val = _RANDOM_554[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_fp_single = _RANDOM_554[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_xcpt_if = _RANDOM_554[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_replay_if = _RANDOM_554[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_555 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_556 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_debug_wdata = {_RANDOM_556[4:0], _RANDOM_555, _RANDOM_554[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_557 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_21_debug_events_fetch_seq = {_RANDOM_557[4:0], _RANDOM_556[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_valid = _RANDOM_557[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_iw_state = _RANDOM_557[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_uopc = _RANDOM_557[16:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_558 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_inst = {_RANDOM_558[16:0], _RANDOM_557[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_559 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_pc = {_RANDOM_559[24:0], _RANDOM_558[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_560 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_fu_code = {_RANDOM_560[0], _RANDOM_559[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_br_type = _RANDOM_560[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_op1_sel = _RANDOM_560[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_op2_sel = _RANDOM_560[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_imm_sel = _RANDOM_560[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_op_fcn = _RANDOM_560[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_fcn_dw = _RANDOM_560[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_rf_wen = _RANDOM_560[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_csr_cmd = _RANDOM_560[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_is_load = _RANDOM_560[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_is_sta = _RANDOM_560[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ctrl_is_std = _RANDOM_560[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_wakeup_delay = _RANDOM_560[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_allocate_brtag = _RANDOM_560[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_br_or_jmp = _RANDOM_560[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_jump = _RANDOM_560[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_jal = _RANDOM_560[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_ret = _RANDOM_560[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_561 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_call = _RANDOM_561[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_mask = _RANDOM_561[8:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_tag = _RANDOM_561[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_prediction_bpd_predict_val = _RANDOM_561[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_prediction_bpd_predict_taken = _RANDOM_561[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_prediction_btb_hit = _RANDOM_561[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_prediction_btb_predicted = _RANDOM_561[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_br_prediction_is_br_or_jalr = _RANDOM_561[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stat_brjmp_mispredicted = _RANDOM_561[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stat_btb_made_pred = _RANDOM_561[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stat_btb_mispredicted = _RANDOM_561[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stat_bpd_made_pred = _RANDOM_561[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stat_bpd_mispredicted = _RANDOM_561[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_fetch_pc_lob = _RANDOM_561[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_562 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_imm_packed = {_RANDOM_562[12:0], _RANDOM_561[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_csr_addr = _RANDOM_562[24:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_rob_idx = _RANDOM_562[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_563 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ldq_idx = {_RANDOM_563[2:0], _RANDOM_562[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stq_idx = _RANDOM_563[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_brob_idx = _RANDOM_563[11:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_pdst = _RANDOM_563[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_pop1 = _RANDOM_563[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_564 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_pop2 = {_RANDOM_564[0], _RANDOM_563[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_pop3 = _RANDOM_564[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_prs1_busy = _RANDOM_564[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_prs2_busy = _RANDOM_564[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_prs3_busy = _RANDOM_564[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_stale_pdst = _RANDOM_564[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_exception = _RANDOM_564[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_565 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_566 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_exc_cause = {_RANDOM_566[18:0], _RANDOM_565, _RANDOM_564[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_bypassable = _RANDOM_566[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_mem_cmd = _RANDOM_566[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_mem_typ = _RANDOM_566[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_fence = _RANDOM_566[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_fencei = _RANDOM_566[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_store = _RANDOM_566[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_amo = _RANDOM_566[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_load = _RANDOM_566[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_567 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_is_unique = _RANDOM_567[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_flush_on_commit = _RANDOM_567[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ldst = _RANDOM_567[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_lrs1 = _RANDOM_567[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_lrs2 = _RANDOM_567[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_lrs3 = _RANDOM_567[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_ldst_val = _RANDOM_567[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_dst_rtype = _RANDOM_567[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_lrs1_rtype = _RANDOM_567[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_568 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_lrs2_rtype = {_RANDOM_568[0], _RANDOM_567[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_frs3_en = _RANDOM_568[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_fp_val = _RANDOM_568[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_fp_single = _RANDOM_568[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_xcpt_if = _RANDOM_568[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_replay_if = _RANDOM_568[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_569 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_570 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_debug_wdata = {_RANDOM_570[5:0], _RANDOM_569, _RANDOM_568[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_571 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_22_debug_events_fetch_seq = {_RANDOM_571[5:0], _RANDOM_570[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_valid = _RANDOM_571[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_iw_state = _RANDOM_571[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_uopc = _RANDOM_571[17:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_572 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_inst = {_RANDOM_572[17:0], _RANDOM_571[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_573 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_pc = {_RANDOM_573[25:0], _RANDOM_572[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_574 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_fu_code = {_RANDOM_574[1:0], _RANDOM_573[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_br_type = _RANDOM_574[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_op1_sel = _RANDOM_574[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_op2_sel = _RANDOM_574[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_imm_sel = _RANDOM_574[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_op_fcn = _RANDOM_574[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_fcn_dw = _RANDOM_574[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_rf_wen = _RANDOM_574[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_csr_cmd = _RANDOM_574[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_is_load = _RANDOM_574[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_is_sta = _RANDOM_574[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ctrl_is_std = _RANDOM_574[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_wakeup_delay = _RANDOM_574[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_allocate_brtag = _RANDOM_574[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_br_or_jmp = _RANDOM_574[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_jump = _RANDOM_574[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_jal = _RANDOM_574[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_575 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_ret = _RANDOM_575[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_call = _RANDOM_575[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_mask = _RANDOM_575[9:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_tag = _RANDOM_575[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_prediction_bpd_predict_val = _RANDOM_575[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_prediction_bpd_predict_taken = _RANDOM_575[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_prediction_btb_hit = _RANDOM_575[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_prediction_btb_predicted = _RANDOM_575[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_br_prediction_is_br_or_jalr = _RANDOM_575[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stat_brjmp_mispredicted = _RANDOM_575[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stat_btb_made_pred = _RANDOM_575[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stat_btb_mispredicted = _RANDOM_575[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stat_bpd_made_pred = _RANDOM_575[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stat_bpd_mispredicted = _RANDOM_575[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_fetch_pc_lob = _RANDOM_575[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_576 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_imm_packed = {_RANDOM_576[13:0], _RANDOM_575[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_csr_addr = _RANDOM_576[25:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_rob_idx = _RANDOM_576[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_577 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ldq_idx = _RANDOM_577[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stq_idx = _RANDOM_577[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_brob_idx = _RANDOM_577[12:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_pdst = _RANDOM_577[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_pop1 = _RANDOM_577[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_578 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_pop2 = {_RANDOM_578[1:0], _RANDOM_577[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_pop3 = _RANDOM_578[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_prs1_busy = _RANDOM_578[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_prs2_busy = _RANDOM_578[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_prs3_busy = _RANDOM_578[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_stale_pdst = _RANDOM_578[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_exception = _RANDOM_578[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_579 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_580 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_exc_cause = {_RANDOM_580[19:0], _RANDOM_579, _RANDOM_578[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_bypassable = _RANDOM_580[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_mem_cmd = _RANDOM_580[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_mem_typ = _RANDOM_580[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_fence = _RANDOM_580[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_fencei = _RANDOM_580[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_store = _RANDOM_580[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_amo = _RANDOM_580[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_581 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_load = _RANDOM_581[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_is_unique = _RANDOM_581[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_flush_on_commit = _RANDOM_581[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ldst = _RANDOM_581[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_lrs1 = _RANDOM_581[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_lrs2 = _RANDOM_581[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_lrs3 = _RANDOM_581[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_ldst_val = _RANDOM_581[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_dst_rtype = _RANDOM_581[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_lrs1_rtype = _RANDOM_581[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_582 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_lrs2_rtype = _RANDOM_582[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_frs3_en = _RANDOM_582[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_fp_val = _RANDOM_582[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_fp_single = _RANDOM_582[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_xcpt_if = _RANDOM_582[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_replay_if = _RANDOM_582[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_583 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_584 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_debug_wdata = {_RANDOM_584[6:0], _RANDOM_583, _RANDOM_582[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        _RANDOM_585 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_26182_23_debug_events_fetch_seq = {_RANDOM_585[6:0], _RANDOM_584[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:189:5
        T_35634_0 = _RANDOM_585[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_1 = _RANDOM_585[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_2 = _RANDOM_585[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_3 = _RANDOM_585[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_4 = _RANDOM_585[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_5 = _RANDOM_585[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_6 = _RANDOM_585[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_7 = _RANDOM_585[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_8 = _RANDOM_585[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_9 = _RANDOM_585[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_10 = _RANDOM_585[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_11 = _RANDOM_585[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_12 = _RANDOM_585[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_13 = _RANDOM_585[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_14 = _RANDOM_585[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_15 = _RANDOM_585[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_16 = _RANDOM_585[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_17 = _RANDOM_585[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_18 = _RANDOM_585[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_19 = _RANDOM_585[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_20 = _RANDOM_585[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_21 = _RANDOM_585[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_22 = _RANDOM_585[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_35634_23 = _RANDOM_585[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1555:5
        T_38110_0_valid = _RANDOM_585[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_586 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_iw_state = _RANDOM_586[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_uopc = _RANDOM_586[10:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_587 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_inst = {_RANDOM_587[10:0], _RANDOM_586[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_588 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_pc = {_RANDOM_588[18:0], _RANDOM_587[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_fu_code = _RANDOM_588[26:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_br_type = _RANDOM_588[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_589 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_op1_sel = {_RANDOM_589[0], _RANDOM_588[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_op2_sel = _RANDOM_589[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_imm_sel = _RANDOM_589[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_op_fcn = _RANDOM_589[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_fcn_dw = _RANDOM_589[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_rf_wen = _RANDOM_589[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_csr_cmd = _RANDOM_589[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_is_load = _RANDOM_589[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_is_sta = _RANDOM_589[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ctrl_is_std = _RANDOM_589[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_wakeup_delay = _RANDOM_589[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_allocate_brtag = _RANDOM_589[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_br_or_jmp = _RANDOM_589[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_jump = _RANDOM_589[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_jal = _RANDOM_589[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_ret = _RANDOM_589[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_call = _RANDOM_589[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_590 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_mask = {_RANDOM_590[2:0], _RANDOM_589[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_tag = _RANDOM_590[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_prediction_bpd_predict_val = _RANDOM_590[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_prediction_bpd_predict_taken = _RANDOM_590[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_prediction_btb_hit = _RANDOM_590[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_prediction_btb_predicted = _RANDOM_590[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_br_prediction_is_br_or_jalr = _RANDOM_590[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stat_brjmp_mispredicted = _RANDOM_590[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stat_btb_made_pred = _RANDOM_590[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stat_btb_mispredicted = _RANDOM_590[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stat_bpd_made_pred = _RANDOM_590[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stat_bpd_mispredicted = _RANDOM_590[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_fetch_pc_lob = _RANDOM_590[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_591 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_imm_packed = {_RANDOM_591[6:0], _RANDOM_590[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_csr_addr = _RANDOM_591[18:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_rob_idx = _RANDOM_591[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ldq_idx = _RANDOM_591[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_592 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stq_idx = {_RANDOM_592[0], _RANDOM_591[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_brob_idx = _RANDOM_592[5:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_pdst = _RANDOM_592[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_pop1 = _RANDOM_592[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_pop2 = _RANDOM_592[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_593 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_pop3 = {_RANDOM_593[1:0], _RANDOM_592[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_prs1_busy = _RANDOM_593[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_prs2_busy = _RANDOM_593[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_prs3_busy = _RANDOM_593[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_stale_pdst = _RANDOM_593[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_exception = _RANDOM_593[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_594 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_595 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_exc_cause = {_RANDOM_595[12:0], _RANDOM_594, _RANDOM_593[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_bypassable = _RANDOM_595[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_mem_cmd = _RANDOM_595[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_mem_typ = _RANDOM_595[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_fence = _RANDOM_595[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_fencei = _RANDOM_595[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_store = _RANDOM_595[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_amo = _RANDOM_595[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_load = _RANDOM_595[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_is_unique = _RANDOM_595[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_flush_on_commit = _RANDOM_595[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_596 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ldst = {_RANDOM_596[1:0], _RANDOM_595[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_lrs1 = _RANDOM_596[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_lrs2 = _RANDOM_596[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_lrs3 = _RANDOM_596[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_ldst_val = _RANDOM_596[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_dst_rtype = _RANDOM_596[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_lrs1_rtype = _RANDOM_596[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_lrs2_rtype = _RANDOM_596[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_frs3_en = _RANDOM_596[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_fp_val = _RANDOM_596[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_fp_single = _RANDOM_596[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_xcpt_if = _RANDOM_596[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_replay_if = _RANDOM_596[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_597 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_598 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_debug_wdata = {_RANDOM_598, _RANDOM_597};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_599 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_0_debug_events_fetch_seq = _RANDOM_599;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_600 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_valid = _RANDOM_600[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_iw_state = _RANDOM_600[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_uopc = _RANDOM_600[11:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_601 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_inst = {_RANDOM_601[11:0], _RANDOM_600[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_602 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_pc = {_RANDOM_602[19:0], _RANDOM_601[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_fu_code = _RANDOM_602[27:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_br_type = _RANDOM_602[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_603 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_op1_sel = _RANDOM_603[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_op2_sel = _RANDOM_603[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_imm_sel = _RANDOM_603[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_op_fcn = _RANDOM_603[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_fcn_dw = _RANDOM_603[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_rf_wen = _RANDOM_603[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_csr_cmd = _RANDOM_603[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_is_load = _RANDOM_603[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_is_sta = _RANDOM_603[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ctrl_is_std = _RANDOM_603[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_wakeup_delay = _RANDOM_603[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_allocate_brtag = _RANDOM_603[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_br_or_jmp = _RANDOM_603[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_jump = _RANDOM_603[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_jal = _RANDOM_603[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_ret = _RANDOM_603[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_call = _RANDOM_603[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_604 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_mask = {_RANDOM_604[3:0], _RANDOM_603[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_tag = _RANDOM_604[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_prediction_bpd_predict_val = _RANDOM_604[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_prediction_bpd_predict_taken = _RANDOM_604[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_prediction_btb_hit = _RANDOM_604[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_prediction_btb_predicted = _RANDOM_604[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_br_prediction_is_br_or_jalr = _RANDOM_604[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stat_brjmp_mispredicted = _RANDOM_604[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stat_btb_made_pred = _RANDOM_604[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stat_btb_mispredicted = _RANDOM_604[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stat_bpd_made_pred = _RANDOM_604[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stat_bpd_mispredicted = _RANDOM_604[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_fetch_pc_lob = _RANDOM_604[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_605 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_imm_packed = {_RANDOM_605[7:0], _RANDOM_604[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_csr_addr = _RANDOM_605[19:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_rob_idx = _RANDOM_605[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ldq_idx = _RANDOM_605[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_606 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stq_idx = {_RANDOM_606[1:0], _RANDOM_605[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_brob_idx = _RANDOM_606[6:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_pdst = _RANDOM_606[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_pop1 = _RANDOM_606[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_pop2 = _RANDOM_606[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_607 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_pop3 = {_RANDOM_607[2:0], _RANDOM_606[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_prs1_busy = _RANDOM_607[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_prs2_busy = _RANDOM_607[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_prs3_busy = _RANDOM_607[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_stale_pdst = _RANDOM_607[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_exception = _RANDOM_607[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_608 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_609 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_exc_cause = {_RANDOM_609[13:0], _RANDOM_608, _RANDOM_607[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_bypassable = _RANDOM_609[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_mem_cmd = _RANDOM_609[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_mem_typ = _RANDOM_609[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_fence = _RANDOM_609[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_fencei = _RANDOM_609[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_store = _RANDOM_609[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_amo = _RANDOM_609[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_load = _RANDOM_609[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_is_unique = _RANDOM_609[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_flush_on_commit = _RANDOM_609[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_610 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ldst = {_RANDOM_610[2:0], _RANDOM_609[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_lrs1 = _RANDOM_610[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_lrs2 = _RANDOM_610[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_lrs3 = _RANDOM_610[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_ldst_val = _RANDOM_610[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_dst_rtype = _RANDOM_610[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_lrs1_rtype = _RANDOM_610[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_lrs2_rtype = _RANDOM_610[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_frs3_en = _RANDOM_610[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_fp_val = _RANDOM_610[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_fp_single = _RANDOM_610[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_xcpt_if = _RANDOM_610[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_611 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_replay_if = _RANDOM_611[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_612 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_613 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_debug_wdata = {_RANDOM_613[0], _RANDOM_612, _RANDOM_611[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_614 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_1_debug_events_fetch_seq = {_RANDOM_614[0], _RANDOM_613[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_valid = _RANDOM_614[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_iw_state = _RANDOM_614[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_uopc = _RANDOM_614[12:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_615 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_inst = {_RANDOM_615[12:0], _RANDOM_614[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_616 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_pc = {_RANDOM_616[20:0], _RANDOM_615[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_fu_code = _RANDOM_616[28:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_617 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_br_type = {_RANDOM_617[0], _RANDOM_616[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_op1_sel = _RANDOM_617[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_op2_sel = _RANDOM_617[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_imm_sel = _RANDOM_617[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_op_fcn = _RANDOM_617[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_fcn_dw = _RANDOM_617[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_rf_wen = _RANDOM_617[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_csr_cmd = _RANDOM_617[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_is_load = _RANDOM_617[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_is_sta = _RANDOM_617[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ctrl_is_std = _RANDOM_617[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_wakeup_delay = _RANDOM_617[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_allocate_brtag = _RANDOM_617[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_br_or_jmp = _RANDOM_617[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_jump = _RANDOM_617[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_jal = _RANDOM_617[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_ret = _RANDOM_617[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_call = _RANDOM_617[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_618 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_mask = {_RANDOM_618[4:0], _RANDOM_617[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_tag = _RANDOM_618[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_prediction_bpd_predict_val = _RANDOM_618[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_prediction_bpd_predict_taken = _RANDOM_618[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_prediction_btb_hit = _RANDOM_618[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_prediction_btb_predicted = _RANDOM_618[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_br_prediction_is_br_or_jalr = _RANDOM_618[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stat_brjmp_mispredicted = _RANDOM_618[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stat_btb_made_pred = _RANDOM_618[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stat_btb_mispredicted = _RANDOM_618[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stat_bpd_made_pred = _RANDOM_618[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stat_bpd_mispredicted = _RANDOM_618[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_fetch_pc_lob = _RANDOM_618[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_619 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_imm_packed = {_RANDOM_619[8:0], _RANDOM_618[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_csr_addr = _RANDOM_619[20:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_rob_idx = _RANDOM_619[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ldq_idx = _RANDOM_619[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_620 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stq_idx = {_RANDOM_620[2:0], _RANDOM_619[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_brob_idx = _RANDOM_620[7:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_pdst = _RANDOM_620[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_pop1 = _RANDOM_620[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_pop2 = _RANDOM_620[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_621 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_pop3 = {_RANDOM_621[3:0], _RANDOM_620[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_prs1_busy = _RANDOM_621[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_prs2_busy = _RANDOM_621[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_prs3_busy = _RANDOM_621[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_stale_pdst = _RANDOM_621[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_exception = _RANDOM_621[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_622 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_623 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_exc_cause = {_RANDOM_623[14:0], _RANDOM_622, _RANDOM_621[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_bypassable = _RANDOM_623[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_mem_cmd = _RANDOM_623[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_mem_typ = _RANDOM_623[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_fence = _RANDOM_623[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_fencei = _RANDOM_623[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_store = _RANDOM_623[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_amo = _RANDOM_623[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_load = _RANDOM_623[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_is_unique = _RANDOM_623[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_flush_on_commit = _RANDOM_623[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_624 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ldst = {_RANDOM_624[3:0], _RANDOM_623[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_lrs1 = _RANDOM_624[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_lrs2 = _RANDOM_624[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_lrs3 = _RANDOM_624[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_ldst_val = _RANDOM_624[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_dst_rtype = _RANDOM_624[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_lrs1_rtype = _RANDOM_624[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_lrs2_rtype = _RANDOM_624[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_frs3_en = _RANDOM_624[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_fp_val = _RANDOM_624[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_fp_single = _RANDOM_624[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_625 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_xcpt_if = _RANDOM_625[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_replay_if = _RANDOM_625[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_626 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_627 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_debug_wdata = {_RANDOM_627[1:0], _RANDOM_626, _RANDOM_625[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_628 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_2_debug_events_fetch_seq = {_RANDOM_628[1:0], _RANDOM_627[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_valid = _RANDOM_628[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_iw_state = _RANDOM_628[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_uopc = _RANDOM_628[13:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_629 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_inst = {_RANDOM_629[13:0], _RANDOM_628[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_630 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_pc = {_RANDOM_630[21:0], _RANDOM_629[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_fu_code = _RANDOM_630[29:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_631 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_br_type = {_RANDOM_631[1:0], _RANDOM_630[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_op1_sel = _RANDOM_631[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_op2_sel = _RANDOM_631[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_imm_sel = _RANDOM_631[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_op_fcn = _RANDOM_631[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_fcn_dw = _RANDOM_631[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_rf_wen = _RANDOM_631[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_csr_cmd = _RANDOM_631[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_is_load = _RANDOM_631[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_is_sta = _RANDOM_631[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ctrl_is_std = _RANDOM_631[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_wakeup_delay = _RANDOM_631[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_allocate_brtag = _RANDOM_631[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_br_or_jmp = _RANDOM_631[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_jump = _RANDOM_631[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_jal = _RANDOM_631[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_ret = _RANDOM_631[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_call = _RANDOM_631[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_632 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_mask = {_RANDOM_632[5:0], _RANDOM_631[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_tag = _RANDOM_632[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_prediction_bpd_predict_val = _RANDOM_632[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_prediction_bpd_predict_taken = _RANDOM_632[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_prediction_btb_hit = _RANDOM_632[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_prediction_btb_predicted = _RANDOM_632[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_br_prediction_is_br_or_jalr = _RANDOM_632[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stat_brjmp_mispredicted = _RANDOM_632[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stat_btb_made_pred = _RANDOM_632[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stat_btb_mispredicted = _RANDOM_632[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stat_bpd_made_pred = _RANDOM_632[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stat_bpd_mispredicted = _RANDOM_632[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_fetch_pc_lob = _RANDOM_632[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_633 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_imm_packed = {_RANDOM_633[9:0], _RANDOM_632[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_csr_addr = _RANDOM_633[21:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_rob_idx = _RANDOM_633[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ldq_idx = _RANDOM_633[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_634 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stq_idx = _RANDOM_634[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_brob_idx = _RANDOM_634[8:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_pdst = _RANDOM_634[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_pop1 = _RANDOM_634[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_pop2 = _RANDOM_634[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_635 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_pop3 = {_RANDOM_635[4:0], _RANDOM_634[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_prs1_busy = _RANDOM_635[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_prs2_busy = _RANDOM_635[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_prs3_busy = _RANDOM_635[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_stale_pdst = _RANDOM_635[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_exception = _RANDOM_635[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_636 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_637 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_exc_cause = {_RANDOM_637[15:0], _RANDOM_636, _RANDOM_635[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_bypassable = _RANDOM_637[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_mem_cmd = _RANDOM_637[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_mem_typ = _RANDOM_637[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_fence = _RANDOM_637[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_fencei = _RANDOM_637[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_store = _RANDOM_637[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_amo = _RANDOM_637[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_load = _RANDOM_637[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_is_unique = _RANDOM_637[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_flush_on_commit = _RANDOM_637[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_638 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ldst = {_RANDOM_638[4:0], _RANDOM_637[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_lrs1 = _RANDOM_638[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_lrs2 = _RANDOM_638[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_lrs3 = _RANDOM_638[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_ldst_val = _RANDOM_638[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_dst_rtype = _RANDOM_638[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_lrs1_rtype = _RANDOM_638[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_lrs2_rtype = _RANDOM_638[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_frs3_en = _RANDOM_638[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_fp_val = _RANDOM_638[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_639 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_fp_single = _RANDOM_639[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_xcpt_if = _RANDOM_639[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_replay_if = _RANDOM_639[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_640 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_641 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_debug_wdata = {_RANDOM_641[2:0], _RANDOM_640, _RANDOM_639[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_642 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_3_debug_events_fetch_seq = {_RANDOM_642[2:0], _RANDOM_641[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_valid = _RANDOM_642[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_iw_state = _RANDOM_642[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_uopc = _RANDOM_642[14:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_643 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_inst = {_RANDOM_643[14:0], _RANDOM_642[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_644 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_pc = {_RANDOM_644[22:0], _RANDOM_643[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_fu_code = _RANDOM_644[30:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_645 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_br_type = {_RANDOM_645[2:0], _RANDOM_644[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_op1_sel = _RANDOM_645[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_op2_sel = _RANDOM_645[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_imm_sel = _RANDOM_645[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_op_fcn = _RANDOM_645[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_fcn_dw = _RANDOM_645[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_rf_wen = _RANDOM_645[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_csr_cmd = _RANDOM_645[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_is_load = _RANDOM_645[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_is_sta = _RANDOM_645[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ctrl_is_std = _RANDOM_645[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_wakeup_delay = _RANDOM_645[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_allocate_brtag = _RANDOM_645[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_br_or_jmp = _RANDOM_645[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_jump = _RANDOM_645[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_jal = _RANDOM_645[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_ret = _RANDOM_645[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_call = _RANDOM_645[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_646 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_mask = {_RANDOM_646[6:0], _RANDOM_645[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_tag = _RANDOM_646[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_prediction_bpd_predict_val = _RANDOM_646[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_prediction_bpd_predict_taken = _RANDOM_646[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_prediction_btb_hit = _RANDOM_646[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_prediction_btb_predicted = _RANDOM_646[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_br_prediction_is_br_or_jalr = _RANDOM_646[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stat_brjmp_mispredicted = _RANDOM_646[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stat_btb_made_pred = _RANDOM_646[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stat_btb_mispredicted = _RANDOM_646[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stat_bpd_made_pred = _RANDOM_646[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stat_bpd_mispredicted = _RANDOM_646[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_fetch_pc_lob = _RANDOM_646[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_647 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_imm_packed = {_RANDOM_647[10:0], _RANDOM_646[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_csr_addr = _RANDOM_647[22:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_rob_idx = _RANDOM_647[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_648 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ldq_idx = {_RANDOM_648[0], _RANDOM_647[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stq_idx = _RANDOM_648[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_brob_idx = _RANDOM_648[9:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_pdst = _RANDOM_648[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_pop1 = _RANDOM_648[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_pop2 = _RANDOM_648[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_649 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_pop3 = {_RANDOM_649[5:0], _RANDOM_648[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_prs1_busy = _RANDOM_649[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_prs2_busy = _RANDOM_649[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_prs3_busy = _RANDOM_649[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_stale_pdst = _RANDOM_649[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_exception = _RANDOM_649[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_650 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_651 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_exc_cause = {_RANDOM_651[16:0], _RANDOM_650, _RANDOM_649[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_bypassable = _RANDOM_651[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_mem_cmd = _RANDOM_651[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_mem_typ = _RANDOM_651[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_fence = _RANDOM_651[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_fencei = _RANDOM_651[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_store = _RANDOM_651[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_amo = _RANDOM_651[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_load = _RANDOM_651[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_is_unique = _RANDOM_651[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_flush_on_commit = _RANDOM_651[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_652 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ldst = _RANDOM_652[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_lrs1 = _RANDOM_652[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_lrs2 = _RANDOM_652[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_lrs3 = _RANDOM_652[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_ldst_val = _RANDOM_652[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_dst_rtype = _RANDOM_652[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_lrs1_rtype = _RANDOM_652[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_lrs2_rtype = _RANDOM_652[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_frs3_en = _RANDOM_652[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_653 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_fp_val = _RANDOM_653[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_fp_single = _RANDOM_653[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_xcpt_if = _RANDOM_653[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_replay_if = _RANDOM_653[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_654 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_655 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_debug_wdata = {_RANDOM_655[3:0], _RANDOM_654, _RANDOM_653[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_656 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_4_debug_events_fetch_seq = {_RANDOM_656[3:0], _RANDOM_655[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_valid = _RANDOM_656[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_iw_state = _RANDOM_656[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_uopc = _RANDOM_656[15:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_657 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_inst = {_RANDOM_657[15:0], _RANDOM_656[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_658 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_pc = {_RANDOM_658[23:0], _RANDOM_657[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_fu_code = _RANDOM_658[31:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_659 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_br_type = _RANDOM_659[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_op1_sel = _RANDOM_659[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_op2_sel = _RANDOM_659[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_imm_sel = _RANDOM_659[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_op_fcn = _RANDOM_659[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_fcn_dw = _RANDOM_659[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_rf_wen = _RANDOM_659[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_csr_cmd = _RANDOM_659[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_is_load = _RANDOM_659[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_is_sta = _RANDOM_659[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ctrl_is_std = _RANDOM_659[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_wakeup_delay = _RANDOM_659[25:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_allocate_brtag = _RANDOM_659[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_br_or_jmp = _RANDOM_659[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_jump = _RANDOM_659[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_jal = _RANDOM_659[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_ret = _RANDOM_659[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_call = _RANDOM_659[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_660 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_mask = _RANDOM_660[7:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_tag = _RANDOM_660[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_prediction_bpd_predict_val = _RANDOM_660[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_prediction_bpd_predict_taken = _RANDOM_660[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_prediction_btb_hit = _RANDOM_660[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_prediction_btb_predicted = _RANDOM_660[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_br_prediction_is_br_or_jalr = _RANDOM_660[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stat_brjmp_mispredicted = _RANDOM_660[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stat_btb_made_pred = _RANDOM_660[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stat_btb_mispredicted = _RANDOM_660[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stat_bpd_made_pred = _RANDOM_660[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stat_bpd_mispredicted = _RANDOM_660[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_fetch_pc_lob = _RANDOM_660[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_661 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_imm_packed = {_RANDOM_661[11:0], _RANDOM_660[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_csr_addr = _RANDOM_661[23:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_rob_idx = _RANDOM_661[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_662 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ldq_idx = {_RANDOM_662[1:0], _RANDOM_661[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stq_idx = _RANDOM_662[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_brob_idx = _RANDOM_662[10:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_pdst = _RANDOM_662[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_pop1 = _RANDOM_662[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_pop2 = _RANDOM_662[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_663 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_pop3 = _RANDOM_663[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_prs1_busy = _RANDOM_663[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_prs2_busy = _RANDOM_663[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_prs3_busy = _RANDOM_663[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_stale_pdst = _RANDOM_663[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_exception = _RANDOM_663[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_664 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_665 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_exc_cause = {_RANDOM_665[17:0], _RANDOM_664, _RANDOM_663[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_bypassable = _RANDOM_665[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_mem_cmd = _RANDOM_665[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_mem_typ = _RANDOM_665[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_fence = _RANDOM_665[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_fencei = _RANDOM_665[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_store = _RANDOM_665[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_amo = _RANDOM_665[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_load = _RANDOM_665[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_is_unique = _RANDOM_665[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_666 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_flush_on_commit = _RANDOM_666[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ldst = _RANDOM_666[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_lrs1 = _RANDOM_666[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_lrs2 = _RANDOM_666[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_lrs3 = _RANDOM_666[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_ldst_val = _RANDOM_666[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_dst_rtype = _RANDOM_666[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_lrs1_rtype = _RANDOM_666[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_lrs2_rtype = _RANDOM_666[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_667 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_frs3_en = _RANDOM_667[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_fp_val = _RANDOM_667[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_fp_single = _RANDOM_667[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_xcpt_if = _RANDOM_667[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_replay_if = _RANDOM_667[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_668 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_669 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_debug_wdata = {_RANDOM_669[4:0], _RANDOM_668, _RANDOM_667[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_670 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_5_debug_events_fetch_seq = {_RANDOM_670[4:0], _RANDOM_669[31:5]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_valid = _RANDOM_670[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_iw_state = _RANDOM_670[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_uopc = _RANDOM_670[16:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_671 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_inst = {_RANDOM_671[16:0], _RANDOM_670[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_672 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_pc = {_RANDOM_672[24:0], _RANDOM_671[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_673 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_fu_code = {_RANDOM_673[0], _RANDOM_672[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_br_type = _RANDOM_673[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_op1_sel = _RANDOM_673[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_op2_sel = _RANDOM_673[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_imm_sel = _RANDOM_673[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_op_fcn = _RANDOM_673[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_fcn_dw = _RANDOM_673[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_rf_wen = _RANDOM_673[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_csr_cmd = _RANDOM_673[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_is_load = _RANDOM_673[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_is_sta = _RANDOM_673[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ctrl_is_std = _RANDOM_673[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_wakeup_delay = _RANDOM_673[26:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_allocate_brtag = _RANDOM_673[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_br_or_jmp = _RANDOM_673[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_jump = _RANDOM_673[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_jal = _RANDOM_673[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_ret = _RANDOM_673[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_674 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_call = _RANDOM_674[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_mask = _RANDOM_674[8:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_tag = _RANDOM_674[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_prediction_bpd_predict_val = _RANDOM_674[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_prediction_bpd_predict_taken = _RANDOM_674[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_prediction_btb_hit = _RANDOM_674[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_prediction_btb_predicted = _RANDOM_674[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_br_prediction_is_br_or_jalr = _RANDOM_674[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stat_brjmp_mispredicted = _RANDOM_674[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stat_btb_made_pred = _RANDOM_674[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stat_btb_mispredicted = _RANDOM_674[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stat_bpd_made_pred = _RANDOM_674[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stat_bpd_mispredicted = _RANDOM_674[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_fetch_pc_lob = _RANDOM_674[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_675 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_imm_packed = {_RANDOM_675[12:0], _RANDOM_674[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_csr_addr = _RANDOM_675[24:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_rob_idx = _RANDOM_675[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_676 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ldq_idx = {_RANDOM_676[2:0], _RANDOM_675[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stq_idx = _RANDOM_676[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_brob_idx = _RANDOM_676[11:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_pdst = _RANDOM_676[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_pop1 = _RANDOM_676[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_677 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_pop2 = {_RANDOM_677[0], _RANDOM_676[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_pop3 = _RANDOM_677[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_prs1_busy = _RANDOM_677[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_prs2_busy = _RANDOM_677[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_prs3_busy = _RANDOM_677[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_stale_pdst = _RANDOM_677[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_exception = _RANDOM_677[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_678 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_679 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_exc_cause = {_RANDOM_679[18:0], _RANDOM_678, _RANDOM_677[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_bypassable = _RANDOM_679[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_mem_cmd = _RANDOM_679[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_mem_typ = _RANDOM_679[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_fence = _RANDOM_679[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_fencei = _RANDOM_679[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_store = _RANDOM_679[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_amo = _RANDOM_679[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_load = _RANDOM_679[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_680 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_is_unique = _RANDOM_680[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_flush_on_commit = _RANDOM_680[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ldst = _RANDOM_680[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_lrs1 = _RANDOM_680[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_lrs2 = _RANDOM_680[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_lrs3 = _RANDOM_680[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_ldst_val = _RANDOM_680[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_dst_rtype = _RANDOM_680[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_lrs1_rtype = _RANDOM_680[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_681 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_lrs2_rtype = {_RANDOM_681[0], _RANDOM_680[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_frs3_en = _RANDOM_681[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_fp_val = _RANDOM_681[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_fp_single = _RANDOM_681[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_xcpt_if = _RANDOM_681[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_replay_if = _RANDOM_681[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_682 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_683 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_debug_wdata = {_RANDOM_683[5:0], _RANDOM_682, _RANDOM_681[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_684 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_6_debug_events_fetch_seq = {_RANDOM_684[5:0], _RANDOM_683[31:6]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_valid = _RANDOM_684[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_iw_state = _RANDOM_684[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_uopc = _RANDOM_684[17:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_685 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_inst = {_RANDOM_685[17:0], _RANDOM_684[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_686 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_pc = {_RANDOM_686[25:0], _RANDOM_685[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_687 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_fu_code = {_RANDOM_687[1:0], _RANDOM_686[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_br_type = _RANDOM_687[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_op1_sel = _RANDOM_687[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_op2_sel = _RANDOM_687[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_imm_sel = _RANDOM_687[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_op_fcn = _RANDOM_687[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_fcn_dw = _RANDOM_687[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_rf_wen = _RANDOM_687[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_csr_cmd = _RANDOM_687[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_is_load = _RANDOM_687[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_is_sta = _RANDOM_687[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ctrl_is_std = _RANDOM_687[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_wakeup_delay = _RANDOM_687[27:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_allocate_brtag = _RANDOM_687[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_br_or_jmp = _RANDOM_687[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_jump = _RANDOM_687[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_jal = _RANDOM_687[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_688 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_ret = _RANDOM_688[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_call = _RANDOM_688[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_mask = _RANDOM_688[9:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_tag = _RANDOM_688[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_prediction_bpd_predict_val = _RANDOM_688[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_prediction_bpd_predict_taken = _RANDOM_688[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_prediction_btb_hit = _RANDOM_688[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_prediction_btb_predicted = _RANDOM_688[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_br_prediction_is_br_or_jalr = _RANDOM_688[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stat_brjmp_mispredicted = _RANDOM_688[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stat_btb_made_pred = _RANDOM_688[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stat_btb_mispredicted = _RANDOM_688[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stat_bpd_made_pred = _RANDOM_688[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stat_bpd_mispredicted = _RANDOM_688[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_fetch_pc_lob = _RANDOM_688[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_689 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_imm_packed = {_RANDOM_689[13:0], _RANDOM_688[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_csr_addr = _RANDOM_689[25:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_rob_idx = _RANDOM_689[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_690 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ldq_idx = _RANDOM_690[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stq_idx = _RANDOM_690[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_brob_idx = _RANDOM_690[12:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_pdst = _RANDOM_690[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_pop1 = _RANDOM_690[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_691 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_pop2 = {_RANDOM_691[1:0], _RANDOM_690[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_pop3 = _RANDOM_691[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_prs1_busy = _RANDOM_691[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_prs2_busy = _RANDOM_691[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_prs3_busy = _RANDOM_691[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_stale_pdst = _RANDOM_691[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_exception = _RANDOM_691[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_692 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_693 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_exc_cause = {_RANDOM_693[19:0], _RANDOM_692, _RANDOM_691[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_bypassable = _RANDOM_693[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_mem_cmd = _RANDOM_693[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_mem_typ = _RANDOM_693[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_fence = _RANDOM_693[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_fencei = _RANDOM_693[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_store = _RANDOM_693[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_amo = _RANDOM_693[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_694 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_load = _RANDOM_694[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_is_unique = _RANDOM_694[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_flush_on_commit = _RANDOM_694[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ldst = _RANDOM_694[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_lrs1 = _RANDOM_694[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_lrs2 = _RANDOM_694[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_lrs3 = _RANDOM_694[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_ldst_val = _RANDOM_694[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_dst_rtype = _RANDOM_694[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_lrs1_rtype = _RANDOM_694[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_695 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_lrs2_rtype = _RANDOM_695[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_frs3_en = _RANDOM_695[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_fp_val = _RANDOM_695[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_fp_single = _RANDOM_695[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_xcpt_if = _RANDOM_695[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_replay_if = _RANDOM_695[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_696 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_697 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_debug_wdata = {_RANDOM_697[6:0], _RANDOM_696, _RANDOM_695[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_698 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_7_debug_events_fetch_seq = {_RANDOM_698[6:0], _RANDOM_697[31:7]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_valid = _RANDOM_698[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_iw_state = _RANDOM_698[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_uopc = _RANDOM_698[18:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_699 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_inst = {_RANDOM_699[18:0], _RANDOM_698[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_700 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_pc = {_RANDOM_700[26:0], _RANDOM_699[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_701 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_fu_code = {_RANDOM_701[2:0], _RANDOM_700[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_br_type = _RANDOM_701[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_op1_sel = _RANDOM_701[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_op2_sel = _RANDOM_701[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_imm_sel = _RANDOM_701[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_op_fcn = _RANDOM_701[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_fcn_dw = _RANDOM_701[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_rf_wen = _RANDOM_701[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_csr_cmd = _RANDOM_701[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_is_load = _RANDOM_701[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_is_sta = _RANDOM_701[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ctrl_is_std = _RANDOM_701[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_wakeup_delay = _RANDOM_701[28:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_allocate_brtag = _RANDOM_701[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_br_or_jmp = _RANDOM_701[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_jump = _RANDOM_701[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_702 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_jal = _RANDOM_702[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_ret = _RANDOM_702[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_call = _RANDOM_702[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_mask = _RANDOM_702[10:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_tag = _RANDOM_702[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_prediction_bpd_predict_val = _RANDOM_702[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_prediction_bpd_predict_taken = _RANDOM_702[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_prediction_btb_hit = _RANDOM_702[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_prediction_btb_predicted = _RANDOM_702[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_br_prediction_is_br_or_jalr = _RANDOM_702[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stat_brjmp_mispredicted = _RANDOM_702[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stat_btb_made_pred = _RANDOM_702[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stat_btb_mispredicted = _RANDOM_702[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stat_bpd_made_pred = _RANDOM_702[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stat_bpd_mispredicted = _RANDOM_702[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_fetch_pc_lob = _RANDOM_702[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_703 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_imm_packed = {_RANDOM_703[14:0], _RANDOM_702[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_csr_addr = _RANDOM_703[26:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_704 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_rob_idx = {_RANDOM_704[0], _RANDOM_703[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ldq_idx = _RANDOM_704[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stq_idx = _RANDOM_704[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_brob_idx = _RANDOM_704[13:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_pdst = _RANDOM_704[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_pop1 = _RANDOM_704[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_705 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_pop2 = {_RANDOM_705[2:0], _RANDOM_704[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_pop3 = _RANDOM_705[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_prs1_busy = _RANDOM_705[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_prs2_busy = _RANDOM_705[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_prs3_busy = _RANDOM_705[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_stale_pdst = _RANDOM_705[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_exception = _RANDOM_705[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_706 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_707 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_exc_cause = {_RANDOM_707[20:0], _RANDOM_706, _RANDOM_705[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_bypassable = _RANDOM_707[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_mem_cmd = _RANDOM_707[25:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_mem_typ = _RANDOM_707[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_fence = _RANDOM_707[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_fencei = _RANDOM_707[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_store = _RANDOM_707[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_708 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_amo = _RANDOM_708[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_load = _RANDOM_708[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_is_unique = _RANDOM_708[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_flush_on_commit = _RANDOM_708[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ldst = _RANDOM_708[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_lrs1 = _RANDOM_708[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_lrs2 = _RANDOM_708[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_lrs3 = _RANDOM_708[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_ldst_val = _RANDOM_708[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_dst_rtype = _RANDOM_708[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_709 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_lrs1_rtype = {_RANDOM_709[0], _RANDOM_708[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_lrs2_rtype = _RANDOM_709[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_frs3_en = _RANDOM_709[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_fp_val = _RANDOM_709[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_fp_single = _RANDOM_709[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_xcpt_if = _RANDOM_709[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_replay_if = _RANDOM_709[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_710 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_711 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_debug_wdata = {_RANDOM_711[7:0], _RANDOM_710, _RANDOM_709[31:8]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_712 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_8_debug_events_fetch_seq = {_RANDOM_712[7:0], _RANDOM_711[31:8]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_valid = _RANDOM_712[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_iw_state = _RANDOM_712[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_uopc = _RANDOM_712[19:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_713 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_inst = {_RANDOM_713[19:0], _RANDOM_712[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_714 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_pc = {_RANDOM_714[27:0], _RANDOM_713[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_715 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_fu_code = {_RANDOM_715[3:0], _RANDOM_714[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_br_type = _RANDOM_715[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_op1_sel = _RANDOM_715[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_op2_sel = _RANDOM_715[12:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_imm_sel = _RANDOM_715[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_op_fcn = _RANDOM_715[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_fcn_dw = _RANDOM_715[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_rf_wen = _RANDOM_715[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_csr_cmd = _RANDOM_715[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_is_load = _RANDOM_715[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_is_sta = _RANDOM_715[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ctrl_is_std = _RANDOM_715[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_wakeup_delay = _RANDOM_715[29:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_allocate_brtag = _RANDOM_715[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_br_or_jmp = _RANDOM_715[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_716 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_jump = _RANDOM_716[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_jal = _RANDOM_716[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_ret = _RANDOM_716[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_call = _RANDOM_716[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_mask = _RANDOM_716[11:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_tag = _RANDOM_716[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_prediction_bpd_predict_val = _RANDOM_716[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_prediction_bpd_predict_taken = _RANDOM_716[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_prediction_btb_hit = _RANDOM_716[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_prediction_btb_predicted = _RANDOM_716[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_br_prediction_is_br_or_jalr = _RANDOM_716[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stat_brjmp_mispredicted = _RANDOM_716[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stat_btb_made_pred = _RANDOM_716[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stat_btb_mispredicted = _RANDOM_716[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stat_bpd_made_pred = _RANDOM_716[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stat_bpd_mispredicted = _RANDOM_716[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_fetch_pc_lob = _RANDOM_716[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_717 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_imm_packed = {_RANDOM_717[15:0], _RANDOM_716[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_csr_addr = _RANDOM_717[27:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_718 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_rob_idx = {_RANDOM_718[1:0], _RANDOM_717[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ldq_idx = _RANDOM_718[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stq_idx = _RANDOM_718[9:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_brob_idx = _RANDOM_718[14:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_pdst = _RANDOM_718[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_pop1 = _RANDOM_718[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_719 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_pop2 = {_RANDOM_719[3:0], _RANDOM_718[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_pop3 = _RANDOM_719[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_prs1_busy = _RANDOM_719[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_prs2_busy = _RANDOM_719[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_prs3_busy = _RANDOM_719[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_stale_pdst = _RANDOM_719[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_exception = _RANDOM_719[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_720 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_721 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_exc_cause = {_RANDOM_721[21:0], _RANDOM_720, _RANDOM_719[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_bypassable = _RANDOM_721[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_mem_cmd = _RANDOM_721[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_mem_typ = _RANDOM_721[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_fence = _RANDOM_721[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_fencei = _RANDOM_721[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_722 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_store = _RANDOM_722[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_amo = _RANDOM_722[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_load = _RANDOM_722[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_is_unique = _RANDOM_722[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_flush_on_commit = _RANDOM_722[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ldst = _RANDOM_722[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_lrs1 = _RANDOM_722[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_lrs2 = _RANDOM_722[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_lrs3 = _RANDOM_722[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_ldst_val = _RANDOM_722[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_dst_rtype = _RANDOM_722[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_723 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_lrs1_rtype = _RANDOM_723[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_lrs2_rtype = _RANDOM_723[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_frs3_en = _RANDOM_723[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_fp_val = _RANDOM_723[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_fp_single = _RANDOM_723[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_xcpt_if = _RANDOM_723[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_replay_if = _RANDOM_723[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_724 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_725 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_debug_wdata = {_RANDOM_725[8:0], _RANDOM_724, _RANDOM_723[31:9]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_726 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_9_debug_events_fetch_seq = {_RANDOM_726[8:0], _RANDOM_725[31:9]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_valid = _RANDOM_726[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_iw_state = _RANDOM_726[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_uopc = _RANDOM_726[20:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_727 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_inst = {_RANDOM_727[20:0], _RANDOM_726[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_728 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_pc = {_RANDOM_728[28:0], _RANDOM_727[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_729 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_fu_code = {_RANDOM_729[4:0], _RANDOM_728[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_br_type = _RANDOM_729[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_op1_sel = _RANDOM_729[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_op2_sel = _RANDOM_729[13:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_imm_sel = _RANDOM_729[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_op_fcn = _RANDOM_729[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_fcn_dw = _RANDOM_729[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_rf_wen = _RANDOM_729[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_csr_cmd = _RANDOM_729[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_is_load = _RANDOM_729[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_is_sta = _RANDOM_729[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ctrl_is_std = _RANDOM_729[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_wakeup_delay = _RANDOM_729[30:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_allocate_brtag = _RANDOM_729[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_730 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_br_or_jmp = _RANDOM_730[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_jump = _RANDOM_730[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_jal = _RANDOM_730[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_ret = _RANDOM_730[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_call = _RANDOM_730[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_mask = _RANDOM_730[12:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_tag = _RANDOM_730[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_prediction_bpd_predict_val = _RANDOM_730[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_prediction_bpd_predict_taken = _RANDOM_730[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_prediction_btb_hit = _RANDOM_730[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_prediction_btb_predicted = _RANDOM_730[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_br_prediction_is_br_or_jalr = _RANDOM_730[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stat_brjmp_mispredicted = _RANDOM_730[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stat_btb_made_pred = _RANDOM_730[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stat_btb_mispredicted = _RANDOM_730[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stat_bpd_made_pred = _RANDOM_730[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stat_bpd_mispredicted = _RANDOM_730[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_fetch_pc_lob = _RANDOM_730[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_731 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_imm_packed = {_RANDOM_731[16:0], _RANDOM_730[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_csr_addr = _RANDOM_731[28:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_732 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_rob_idx = {_RANDOM_732[2:0], _RANDOM_731[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ldq_idx = _RANDOM_732[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stq_idx = _RANDOM_732[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_brob_idx = _RANDOM_732[15:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_pdst = _RANDOM_732[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_pop1 = _RANDOM_732[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_733 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_pop2 = {_RANDOM_733[4:0], _RANDOM_732[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_pop3 = _RANDOM_733[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_prs1_busy = _RANDOM_733[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_prs2_busy = _RANDOM_733[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_prs3_busy = _RANDOM_733[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_stale_pdst = _RANDOM_733[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_exception = _RANDOM_733[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_734 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_735 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_exc_cause = {_RANDOM_735[22:0], _RANDOM_734, _RANDOM_733[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_bypassable = _RANDOM_735[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_mem_cmd = _RANDOM_735[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_mem_typ = _RANDOM_735[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_fence = _RANDOM_735[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_736 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_fencei = _RANDOM_736[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_store = _RANDOM_736[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_amo = _RANDOM_736[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_load = _RANDOM_736[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_is_unique = _RANDOM_736[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_flush_on_commit = _RANDOM_736[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ldst = _RANDOM_736[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_lrs1 = _RANDOM_736[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_lrs2 = _RANDOM_736[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_lrs3 = _RANDOM_736[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_ldst_val = _RANDOM_736[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_737 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_dst_rtype = {_RANDOM_737[0], _RANDOM_736[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_lrs1_rtype = _RANDOM_737[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_lrs2_rtype = _RANDOM_737[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_frs3_en = _RANDOM_737[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_fp_val = _RANDOM_737[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_fp_single = _RANDOM_737[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_xcpt_if = _RANDOM_737[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_replay_if = _RANDOM_737[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_738 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_739 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_debug_wdata = {_RANDOM_739[9:0], _RANDOM_738, _RANDOM_737[31:10]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_740 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_10_debug_events_fetch_seq = {_RANDOM_740[9:0], _RANDOM_739[31:10]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_valid = _RANDOM_740[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_iw_state = _RANDOM_740[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_uopc = _RANDOM_740[21:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_741 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_inst = {_RANDOM_741[21:0], _RANDOM_740[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_742 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_pc = {_RANDOM_742[29:0], _RANDOM_741[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_743 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_fu_code = {_RANDOM_743[5:0], _RANDOM_742[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_br_type = _RANDOM_743[9:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_op1_sel = _RANDOM_743[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_op2_sel = _RANDOM_743[14:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_imm_sel = _RANDOM_743[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_op_fcn = _RANDOM_743[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_fcn_dw = _RANDOM_743[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_rf_wen = _RANDOM_743[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_csr_cmd = _RANDOM_743[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_is_load = _RANDOM_743[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_is_sta = _RANDOM_743[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ctrl_is_std = _RANDOM_743[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_wakeup_delay = _RANDOM_743[31:30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_744 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_allocate_brtag = _RANDOM_744[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_br_or_jmp = _RANDOM_744[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_jump = _RANDOM_744[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_jal = _RANDOM_744[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_ret = _RANDOM_744[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_call = _RANDOM_744[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_mask = _RANDOM_744[13:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_tag = _RANDOM_744[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_prediction_bpd_predict_val = _RANDOM_744[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_prediction_bpd_predict_taken = _RANDOM_744[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_prediction_btb_hit = _RANDOM_744[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_prediction_btb_predicted = _RANDOM_744[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_br_prediction_is_br_or_jalr = _RANDOM_744[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stat_brjmp_mispredicted = _RANDOM_744[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stat_btb_made_pred = _RANDOM_744[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stat_btb_mispredicted = _RANDOM_744[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stat_bpd_made_pred = _RANDOM_744[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stat_bpd_mispredicted = _RANDOM_744[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_fetch_pc_lob = _RANDOM_744[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_745 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_imm_packed = {_RANDOM_745[17:0], _RANDOM_744[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_csr_addr = _RANDOM_745[29:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_746 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_rob_idx = {_RANDOM_746[3:0], _RANDOM_745[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ldq_idx = _RANDOM_746[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stq_idx = _RANDOM_746[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_brob_idx = _RANDOM_746[16:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_pdst = _RANDOM_746[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_pop1 = _RANDOM_746[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_747 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_pop2 = {_RANDOM_747[5:0], _RANDOM_746[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_pop3 = _RANDOM_747[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_prs1_busy = _RANDOM_747[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_prs2_busy = _RANDOM_747[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_prs3_busy = _RANDOM_747[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_stale_pdst = _RANDOM_747[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_exception = _RANDOM_747[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_748 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_749 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_exc_cause = {_RANDOM_749[23:0], _RANDOM_748, _RANDOM_747[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_bypassable = _RANDOM_749[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_mem_cmd = _RANDOM_749[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_mem_typ = _RANDOM_749[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_750 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_fence = _RANDOM_750[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_fencei = _RANDOM_750[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_store = _RANDOM_750[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_amo = _RANDOM_750[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_load = _RANDOM_750[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_is_unique = _RANDOM_750[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_flush_on_commit = _RANDOM_750[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ldst = _RANDOM_750[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_lrs1 = _RANDOM_750[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_lrs2 = _RANDOM_750[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_lrs3 = _RANDOM_750[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_ldst_val = _RANDOM_750[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_751 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_dst_rtype = _RANDOM_751[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_lrs1_rtype = _RANDOM_751[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_lrs2_rtype = _RANDOM_751[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_frs3_en = _RANDOM_751[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_fp_val = _RANDOM_751[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_fp_single = _RANDOM_751[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_xcpt_if = _RANDOM_751[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_replay_if = _RANDOM_751[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_752 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_753 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_debug_wdata = {_RANDOM_753[10:0], _RANDOM_752, _RANDOM_751[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_754 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_11_debug_events_fetch_seq = {_RANDOM_754[10:0], _RANDOM_753[31:11]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_valid = _RANDOM_754[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_iw_state = _RANDOM_754[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_uopc = _RANDOM_754[22:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_755 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_inst = {_RANDOM_755[22:0], _RANDOM_754[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_756 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_pc = {_RANDOM_756[30:0], _RANDOM_755[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_757 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_fu_code = {_RANDOM_757[6:0], _RANDOM_756[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_br_type = _RANDOM_757[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_op1_sel = _RANDOM_757[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_op2_sel = _RANDOM_757[15:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_imm_sel = _RANDOM_757[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_op_fcn = _RANDOM_757[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_fcn_dw = _RANDOM_757[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_rf_wen = _RANDOM_757[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_csr_cmd = _RANDOM_757[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_is_load = _RANDOM_757[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_is_sta = _RANDOM_757[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ctrl_is_std = _RANDOM_757[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_758 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_wakeup_delay = {_RANDOM_758[0], _RANDOM_757[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_allocate_brtag = _RANDOM_758[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_br_or_jmp = _RANDOM_758[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_jump = _RANDOM_758[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_jal = _RANDOM_758[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_ret = _RANDOM_758[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_call = _RANDOM_758[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_mask = _RANDOM_758[14:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_tag = _RANDOM_758[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_prediction_bpd_predict_val = _RANDOM_758[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_prediction_bpd_predict_taken = _RANDOM_758[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_prediction_btb_hit = _RANDOM_758[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_prediction_btb_predicted = _RANDOM_758[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_br_prediction_is_br_or_jalr = _RANDOM_758[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stat_brjmp_mispredicted = _RANDOM_758[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stat_btb_made_pred = _RANDOM_758[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stat_btb_mispredicted = _RANDOM_758[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stat_bpd_made_pred = _RANDOM_758[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stat_bpd_mispredicted = _RANDOM_758[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_fetch_pc_lob = _RANDOM_758[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_759 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_imm_packed = {_RANDOM_759[18:0], _RANDOM_758[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_csr_addr = _RANDOM_759[30:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_760 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_rob_idx = {_RANDOM_760[4:0], _RANDOM_759[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ldq_idx = _RANDOM_760[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stq_idx = _RANDOM_760[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_brob_idx = _RANDOM_760[17:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_pdst = _RANDOM_760[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_pop1 = _RANDOM_760[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_761 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_pop2 = _RANDOM_761[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_pop3 = _RANDOM_761[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_prs1_busy = _RANDOM_761[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_prs2_busy = _RANDOM_761[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_prs3_busy = _RANDOM_761[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_stale_pdst = _RANDOM_761[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_exception = _RANDOM_761[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_762 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_763 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_exc_cause = {_RANDOM_763[24:0], _RANDOM_762, _RANDOM_761[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_bypassable = _RANDOM_763[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_mem_cmd = _RANDOM_763[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_764 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_mem_typ = {_RANDOM_764[0], _RANDOM_763[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_fence = _RANDOM_764[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_fencei = _RANDOM_764[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_store = _RANDOM_764[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_amo = _RANDOM_764[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_load = _RANDOM_764[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_is_unique = _RANDOM_764[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_flush_on_commit = _RANDOM_764[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ldst = _RANDOM_764[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_lrs1 = _RANDOM_764[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_lrs2 = _RANDOM_764[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_lrs3 = _RANDOM_764[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_765 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_ldst_val = _RANDOM_765[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_dst_rtype = _RANDOM_765[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_lrs1_rtype = _RANDOM_765[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_lrs2_rtype = _RANDOM_765[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_frs3_en = _RANDOM_765[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_fp_val = _RANDOM_765[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_fp_single = _RANDOM_765[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_xcpt_if = _RANDOM_765[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_replay_if = _RANDOM_765[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_766 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_767 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_debug_wdata = {_RANDOM_767[11:0], _RANDOM_766, _RANDOM_765[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_768 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_12_debug_events_fetch_seq = {_RANDOM_768[11:0], _RANDOM_767[31:12]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_valid = _RANDOM_768[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_iw_state = _RANDOM_768[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_uopc = _RANDOM_768[23:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_769 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_inst = {_RANDOM_769[23:0], _RANDOM_768[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_770 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_pc = {_RANDOM_770, _RANDOM_769[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_771 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_fu_code = _RANDOM_771[7:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_br_type = _RANDOM_771[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_op1_sel = _RANDOM_771[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_op2_sel = _RANDOM_771[16:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_imm_sel = _RANDOM_771[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_op_fcn = _RANDOM_771[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_fcn_dw = _RANDOM_771[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_rf_wen = _RANDOM_771[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_csr_cmd = _RANDOM_771[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_is_load = _RANDOM_771[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_is_sta = _RANDOM_771[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ctrl_is_std = _RANDOM_771[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_772 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_wakeup_delay = _RANDOM_772[1:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_allocate_brtag = _RANDOM_772[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_br_or_jmp = _RANDOM_772[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_jump = _RANDOM_772[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_jal = _RANDOM_772[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_ret = _RANDOM_772[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_call = _RANDOM_772[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_mask = _RANDOM_772[15:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_tag = _RANDOM_772[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_prediction_bpd_predict_val = _RANDOM_772[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_prediction_bpd_predict_taken = _RANDOM_772[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_prediction_btb_hit = _RANDOM_772[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_prediction_btb_predicted = _RANDOM_772[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_br_prediction_is_br_or_jalr = _RANDOM_772[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stat_brjmp_mispredicted = _RANDOM_772[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stat_btb_made_pred = _RANDOM_772[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stat_btb_mispredicted = _RANDOM_772[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stat_bpd_made_pred = _RANDOM_772[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stat_bpd_mispredicted = _RANDOM_772[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_fetch_pc_lob = _RANDOM_772[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_773 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_imm_packed = _RANDOM_773[19:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_csr_addr = _RANDOM_773[31:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_774 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_rob_idx = _RANDOM_774[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ldq_idx = _RANDOM_774[9:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stq_idx = _RANDOM_774[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_brob_idx = _RANDOM_774[18:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_pdst = _RANDOM_774[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_775 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_pop1 = {_RANDOM_775[0], _RANDOM_774[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_pop2 = _RANDOM_775[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_pop3 = _RANDOM_775[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_prs1_busy = _RANDOM_775[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_prs2_busy = _RANDOM_775[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_prs3_busy = _RANDOM_775[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_stale_pdst = _RANDOM_775[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_exception = _RANDOM_775[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_776 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_777 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_exc_cause = {_RANDOM_777[25:0], _RANDOM_776, _RANDOM_775[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_bypassable = _RANDOM_777[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_mem_cmd = _RANDOM_777[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_778 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_mem_typ = {_RANDOM_778[1:0], _RANDOM_777[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_fence = _RANDOM_778[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_fencei = _RANDOM_778[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_store = _RANDOM_778[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_amo = _RANDOM_778[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_load = _RANDOM_778[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_is_unique = _RANDOM_778[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_flush_on_commit = _RANDOM_778[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ldst = _RANDOM_778[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_lrs1 = _RANDOM_778[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_lrs2 = _RANDOM_778[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_779 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_lrs3 = {_RANDOM_779[0], _RANDOM_778[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_ldst_val = _RANDOM_779[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_dst_rtype = _RANDOM_779[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_lrs1_rtype = _RANDOM_779[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_lrs2_rtype = _RANDOM_779[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_frs3_en = _RANDOM_779[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_fp_val = _RANDOM_779[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_fp_single = _RANDOM_779[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_xcpt_if = _RANDOM_779[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_replay_if = _RANDOM_779[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_780 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_781 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_debug_wdata = {_RANDOM_781[12:0], _RANDOM_780, _RANDOM_779[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_782 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_13_debug_events_fetch_seq = {_RANDOM_782[12:0], _RANDOM_781[31:13]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_valid = _RANDOM_782[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_iw_state = _RANDOM_782[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_uopc = _RANDOM_782[24:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_783 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_inst = {_RANDOM_783[24:0], _RANDOM_782[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_784 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_785 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_pc = {_RANDOM_785[0], _RANDOM_784, _RANDOM_783[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_fu_code = _RANDOM_785[8:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_br_type = _RANDOM_785[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_op1_sel = _RANDOM_785[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_op2_sel = _RANDOM_785[17:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_imm_sel = _RANDOM_785[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_op_fcn = _RANDOM_785[24:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_fcn_dw = _RANDOM_785[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_rf_wen = _RANDOM_785[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_csr_cmd = _RANDOM_785[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_is_load = _RANDOM_785[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_is_sta = _RANDOM_785[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_786 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ctrl_is_std = _RANDOM_786[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_wakeup_delay = _RANDOM_786[2:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_allocate_brtag = _RANDOM_786[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_br_or_jmp = _RANDOM_786[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_jump = _RANDOM_786[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_jal = _RANDOM_786[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_ret = _RANDOM_786[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_call = _RANDOM_786[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_mask = _RANDOM_786[16:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_tag = _RANDOM_786[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_prediction_bpd_predict_val = _RANDOM_786[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_prediction_bpd_predict_taken = _RANDOM_786[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_prediction_btb_hit = _RANDOM_786[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_prediction_btb_predicted = _RANDOM_786[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_br_prediction_is_br_or_jalr = _RANDOM_786[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stat_brjmp_mispredicted = _RANDOM_786[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stat_btb_made_pred = _RANDOM_786[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stat_btb_mispredicted = _RANDOM_786[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stat_bpd_made_pred = _RANDOM_786[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stat_bpd_mispredicted = _RANDOM_786[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_787 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_fetch_pc_lob = {_RANDOM_787[0], _RANDOM_786[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_imm_packed = _RANDOM_787[20:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_788 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_csr_addr = {_RANDOM_788[0], _RANDOM_787[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_rob_idx = _RANDOM_788[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ldq_idx = _RANDOM_788[10:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stq_idx = _RANDOM_788[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_brob_idx = _RANDOM_788[19:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_pdst = _RANDOM_788[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_789 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_pop1 = {_RANDOM_789[1:0], _RANDOM_788[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_pop2 = _RANDOM_789[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_pop3 = _RANDOM_789[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_prs1_busy = _RANDOM_789[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_prs2_busy = _RANDOM_789[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_prs3_busy = _RANDOM_789[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_stale_pdst = _RANDOM_789[25:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_exception = _RANDOM_789[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_790 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_791 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_exc_cause = {_RANDOM_791[26:0], _RANDOM_790, _RANDOM_789[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_bypassable = _RANDOM_791[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_mem_cmd = _RANDOM_791[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_792 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_mem_typ = _RANDOM_792[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_fence = _RANDOM_792[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_fencei = _RANDOM_792[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_store = _RANDOM_792[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_amo = _RANDOM_792[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_load = _RANDOM_792[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_is_unique = _RANDOM_792[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_flush_on_commit = _RANDOM_792[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ldst = _RANDOM_792[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_lrs1 = _RANDOM_792[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_lrs2 = _RANDOM_792[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_793 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_lrs3 = {_RANDOM_793[1:0], _RANDOM_792[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_ldst_val = _RANDOM_793[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_dst_rtype = _RANDOM_793[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_lrs1_rtype = _RANDOM_793[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_lrs2_rtype = _RANDOM_793[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_frs3_en = _RANDOM_793[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_fp_val = _RANDOM_793[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_fp_single = _RANDOM_793[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_xcpt_if = _RANDOM_793[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_replay_if = _RANDOM_793[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_794 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_795 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_debug_wdata = {_RANDOM_795[13:0], _RANDOM_794, _RANDOM_793[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_796 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_14_debug_events_fetch_seq = {_RANDOM_796[13:0], _RANDOM_795[31:14]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_valid = _RANDOM_796[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_iw_state = _RANDOM_796[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_uopc = _RANDOM_796[25:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_797 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_inst = {_RANDOM_797[25:0], _RANDOM_796[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_798 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_799 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_pc = {_RANDOM_799[1:0], _RANDOM_798, _RANDOM_797[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_fu_code = _RANDOM_799[9:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_br_type = _RANDOM_799[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_op1_sel = _RANDOM_799[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_op2_sel = _RANDOM_799[18:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_imm_sel = _RANDOM_799[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_op_fcn = _RANDOM_799[25:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_fcn_dw = _RANDOM_799[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_rf_wen = _RANDOM_799[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_csr_cmd = _RANDOM_799[30:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_is_load = _RANDOM_799[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_800 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_is_sta = _RANDOM_800[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ctrl_is_std = _RANDOM_800[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_wakeup_delay = _RANDOM_800[3:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_allocate_brtag = _RANDOM_800[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_br_or_jmp = _RANDOM_800[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_jump = _RANDOM_800[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_jal = _RANDOM_800[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_ret = _RANDOM_800[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_call = _RANDOM_800[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_mask = _RANDOM_800[17:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_tag = _RANDOM_800[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_prediction_bpd_predict_val = _RANDOM_800[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_prediction_bpd_predict_taken = _RANDOM_800[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_prediction_btb_hit = _RANDOM_800[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_prediction_btb_predicted = _RANDOM_800[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_br_prediction_is_br_or_jalr = _RANDOM_800[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stat_brjmp_mispredicted = _RANDOM_800[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stat_btb_made_pred = _RANDOM_800[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stat_btb_mispredicted = _RANDOM_800[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stat_bpd_made_pred = _RANDOM_800[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stat_bpd_mispredicted = _RANDOM_800[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_801 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_fetch_pc_lob = {_RANDOM_801[1:0], _RANDOM_800[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_imm_packed = _RANDOM_801[21:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_802 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_csr_addr = {_RANDOM_802[1:0], _RANDOM_801[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_rob_idx = _RANDOM_802[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ldq_idx = _RANDOM_802[11:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stq_idx = _RANDOM_802[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_brob_idx = _RANDOM_802[20:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_pdst = _RANDOM_802[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_803 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_pop1 = {_RANDOM_803[2:0], _RANDOM_802[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_pop2 = _RANDOM_803[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_pop3 = _RANDOM_803[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_prs1_busy = _RANDOM_803[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_prs2_busy = _RANDOM_803[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_prs3_busy = _RANDOM_803[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_stale_pdst = _RANDOM_803[26:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_exception = _RANDOM_803[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_804 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_805 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_exc_cause = {_RANDOM_805[27:0], _RANDOM_804, _RANDOM_803[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_bypassable = _RANDOM_805[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_806 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_mem_cmd = {_RANDOM_806[0], _RANDOM_805[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_mem_typ = _RANDOM_806[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_fence = _RANDOM_806[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_fencei = _RANDOM_806[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_store = _RANDOM_806[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_amo = _RANDOM_806[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_load = _RANDOM_806[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_is_unique = _RANDOM_806[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_flush_on_commit = _RANDOM_806[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ldst = _RANDOM_806[16:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_lrs1 = _RANDOM_806[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_lrs2 = _RANDOM_806[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_807 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_lrs3 = {_RANDOM_807[2:0], _RANDOM_806[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_ldst_val = _RANDOM_807[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_dst_rtype = _RANDOM_807[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_lrs1_rtype = _RANDOM_807[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_lrs2_rtype = _RANDOM_807[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_frs3_en = _RANDOM_807[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_fp_val = _RANDOM_807[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_fp_single = _RANDOM_807[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_xcpt_if = _RANDOM_807[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_replay_if = _RANDOM_807[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_808 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_809 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_debug_wdata = {_RANDOM_809[14:0], _RANDOM_808, _RANDOM_807[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_810 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_15_debug_events_fetch_seq = {_RANDOM_810[14:0], _RANDOM_809[31:15]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_valid = _RANDOM_810[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_iw_state = _RANDOM_810[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_uopc = _RANDOM_810[26:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_811 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_inst = {_RANDOM_811[26:0], _RANDOM_810[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_812 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_813 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_pc = {_RANDOM_813[2:0], _RANDOM_812, _RANDOM_811[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_fu_code = _RANDOM_813[10:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_br_type = _RANDOM_813[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_op1_sel = _RANDOM_813[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_op2_sel = _RANDOM_813[19:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_imm_sel = _RANDOM_813[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_op_fcn = _RANDOM_813[26:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_fcn_dw = _RANDOM_813[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_rf_wen = _RANDOM_813[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_csr_cmd = _RANDOM_813[31:29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_814 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_is_load = _RANDOM_814[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_is_sta = _RANDOM_814[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ctrl_is_std = _RANDOM_814[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_wakeup_delay = _RANDOM_814[4:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_allocate_brtag = _RANDOM_814[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_br_or_jmp = _RANDOM_814[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_jump = _RANDOM_814[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_jal = _RANDOM_814[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_ret = _RANDOM_814[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_call = _RANDOM_814[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_mask = _RANDOM_814[18:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_tag = _RANDOM_814[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_prediction_bpd_predict_val = _RANDOM_814[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_prediction_bpd_predict_taken = _RANDOM_814[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_prediction_btb_hit = _RANDOM_814[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_prediction_btb_predicted = _RANDOM_814[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_br_prediction_is_br_or_jalr = _RANDOM_814[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stat_brjmp_mispredicted = _RANDOM_814[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stat_btb_made_pred = _RANDOM_814[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stat_btb_mispredicted = _RANDOM_814[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stat_bpd_made_pred = _RANDOM_814[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stat_bpd_mispredicted = _RANDOM_814[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_815 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_fetch_pc_lob = _RANDOM_815[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_imm_packed = _RANDOM_815[22:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_816 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_csr_addr = {_RANDOM_816[2:0], _RANDOM_815[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_rob_idx = _RANDOM_816[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ldq_idx = _RANDOM_816[12:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stq_idx = _RANDOM_816[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_brob_idx = _RANDOM_816[21:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_pdst = _RANDOM_816[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_817 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_pop1 = {_RANDOM_817[3:0], _RANDOM_816[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_pop2 = _RANDOM_817[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_pop3 = _RANDOM_817[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_prs1_busy = _RANDOM_817[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_prs2_busy = _RANDOM_817[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_prs3_busy = _RANDOM_817[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_stale_pdst = _RANDOM_817[27:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_exception = _RANDOM_817[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_818 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_819 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_exc_cause = {_RANDOM_819[28:0], _RANDOM_818, _RANDOM_817[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_bypassable = _RANDOM_819[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_820 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_mem_cmd = {_RANDOM_820[1:0], _RANDOM_819[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_mem_typ = _RANDOM_820[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_fence = _RANDOM_820[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_fencei = _RANDOM_820[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_store = _RANDOM_820[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_amo = _RANDOM_820[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_load = _RANDOM_820[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_is_unique = _RANDOM_820[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_flush_on_commit = _RANDOM_820[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ldst = _RANDOM_820[17:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_lrs1 = _RANDOM_820[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_lrs2 = _RANDOM_820[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_821 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_lrs3 = {_RANDOM_821[3:0], _RANDOM_820[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_ldst_val = _RANDOM_821[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_dst_rtype = _RANDOM_821[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_lrs1_rtype = _RANDOM_821[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_lrs2_rtype = _RANDOM_821[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_frs3_en = _RANDOM_821[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_fp_val = _RANDOM_821[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_fp_single = _RANDOM_821[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_xcpt_if = _RANDOM_821[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_replay_if = _RANDOM_821[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_822 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_823 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_debug_wdata = {_RANDOM_823[15:0], _RANDOM_822, _RANDOM_821[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_824 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_16_debug_events_fetch_seq = {_RANDOM_824[15:0], _RANDOM_823[31:16]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_valid = _RANDOM_824[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_iw_state = _RANDOM_824[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_uopc = _RANDOM_824[27:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_825 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_inst = {_RANDOM_825[27:0], _RANDOM_824[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_826 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_827 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_pc = {_RANDOM_827[3:0], _RANDOM_826, _RANDOM_825[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_fu_code = _RANDOM_827[11:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_br_type = _RANDOM_827[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_op1_sel = _RANDOM_827[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_op2_sel = _RANDOM_827[20:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_imm_sel = _RANDOM_827[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_op_fcn = _RANDOM_827[27:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_fcn_dw = _RANDOM_827[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_rf_wen = _RANDOM_827[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_828 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_csr_cmd = {_RANDOM_828[0], _RANDOM_827[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_is_load = _RANDOM_828[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_is_sta = _RANDOM_828[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ctrl_is_std = _RANDOM_828[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_wakeup_delay = _RANDOM_828[5:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_allocate_brtag = _RANDOM_828[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_br_or_jmp = _RANDOM_828[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_jump = _RANDOM_828[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_jal = _RANDOM_828[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_ret = _RANDOM_828[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_call = _RANDOM_828[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_mask = _RANDOM_828[19:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_tag = _RANDOM_828[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_prediction_bpd_predict_val = _RANDOM_828[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_prediction_bpd_predict_taken = _RANDOM_828[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_prediction_btb_hit = _RANDOM_828[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_prediction_btb_predicted = _RANDOM_828[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_br_prediction_is_br_or_jalr = _RANDOM_828[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stat_brjmp_mispredicted = _RANDOM_828[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stat_btb_made_pred = _RANDOM_828[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stat_btb_mispredicted = _RANDOM_828[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stat_bpd_made_pred = _RANDOM_828[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_829 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stat_bpd_mispredicted = _RANDOM_829[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_fetch_pc_lob = _RANDOM_829[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_imm_packed = _RANDOM_829[23:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_830 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_csr_addr = {_RANDOM_830[3:0], _RANDOM_829[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_rob_idx = _RANDOM_830[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ldq_idx = _RANDOM_830[13:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stq_idx = _RANDOM_830[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_brob_idx = _RANDOM_830[22:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_pdst = _RANDOM_830[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_831 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_pop1 = {_RANDOM_831[4:0], _RANDOM_830[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_pop2 = _RANDOM_831[11:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_pop3 = _RANDOM_831[18:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_prs1_busy = _RANDOM_831[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_prs2_busy = _RANDOM_831[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_prs3_busy = _RANDOM_831[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_stale_pdst = _RANDOM_831[28:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_exception = _RANDOM_831[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_832 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_833 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_exc_cause = {_RANDOM_833[29:0], _RANDOM_832, _RANDOM_831[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_bypassable = _RANDOM_833[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_834 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_mem_cmd = {_RANDOM_834[2:0], _RANDOM_833[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_mem_typ = _RANDOM_834[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_fence = _RANDOM_834[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_fencei = _RANDOM_834[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_store = _RANDOM_834[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_amo = _RANDOM_834[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_load = _RANDOM_834[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_is_unique = _RANDOM_834[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_flush_on_commit = _RANDOM_834[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ldst = _RANDOM_834[18:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_lrs1 = _RANDOM_834[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_lrs2 = _RANDOM_834[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_835 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_lrs3 = {_RANDOM_835[4:0], _RANDOM_834[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_ldst_val = _RANDOM_835[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_dst_rtype = _RANDOM_835[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_lrs1_rtype = _RANDOM_835[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_lrs2_rtype = _RANDOM_835[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_frs3_en = _RANDOM_835[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_fp_val = _RANDOM_835[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_fp_single = _RANDOM_835[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_xcpt_if = _RANDOM_835[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_replay_if = _RANDOM_835[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_836 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_837 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_debug_wdata = {_RANDOM_837[16:0], _RANDOM_836, _RANDOM_835[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_838 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_17_debug_events_fetch_seq = {_RANDOM_838[16:0], _RANDOM_837[31:17]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_valid = _RANDOM_838[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_iw_state = _RANDOM_838[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_uopc = _RANDOM_838[28:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_839 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_inst = {_RANDOM_839[28:0], _RANDOM_838[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_840 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_841 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_pc = {_RANDOM_841[4:0], _RANDOM_840, _RANDOM_839[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_fu_code = _RANDOM_841[12:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_br_type = _RANDOM_841[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_op1_sel = _RANDOM_841[18:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_op2_sel = _RANDOM_841[21:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_imm_sel = _RANDOM_841[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_op_fcn = _RANDOM_841[28:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_fcn_dw = _RANDOM_841[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_rf_wen = _RANDOM_841[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_842 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_csr_cmd = {_RANDOM_842[1:0], _RANDOM_841[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_is_load = _RANDOM_842[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_is_sta = _RANDOM_842[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ctrl_is_std = _RANDOM_842[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_wakeup_delay = _RANDOM_842[6:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_allocate_brtag = _RANDOM_842[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_br_or_jmp = _RANDOM_842[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_jump = _RANDOM_842[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_jal = _RANDOM_842[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_ret = _RANDOM_842[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_call = _RANDOM_842[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_mask = _RANDOM_842[20:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_tag = _RANDOM_842[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_prediction_bpd_predict_val = _RANDOM_842[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_prediction_bpd_predict_taken = _RANDOM_842[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_prediction_btb_hit = _RANDOM_842[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_prediction_btb_predicted = _RANDOM_842[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_br_prediction_is_br_or_jalr = _RANDOM_842[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stat_brjmp_mispredicted = _RANDOM_842[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stat_btb_made_pred = _RANDOM_842[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stat_btb_mispredicted = _RANDOM_842[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_843 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stat_bpd_made_pred = _RANDOM_843[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stat_bpd_mispredicted = _RANDOM_843[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_fetch_pc_lob = _RANDOM_843[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_imm_packed = _RANDOM_843[24:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_844 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_csr_addr = {_RANDOM_844[4:0], _RANDOM_843[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_rob_idx = _RANDOM_844[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ldq_idx = _RANDOM_844[14:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stq_idx = _RANDOM_844[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_brob_idx = _RANDOM_844[23:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_pdst = _RANDOM_844[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_845 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_pop1 = {_RANDOM_845[5:0], _RANDOM_844[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_pop2 = _RANDOM_845[12:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_pop3 = _RANDOM_845[19:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_prs1_busy = _RANDOM_845[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_prs2_busy = _RANDOM_845[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_prs3_busy = _RANDOM_845[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_stale_pdst = _RANDOM_845[29:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_exception = _RANDOM_845[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_846 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_847 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_exc_cause = {_RANDOM_847[30:0], _RANDOM_846, _RANDOM_845[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_bypassable = _RANDOM_847[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_848 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_mem_cmd = _RANDOM_848[3:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_mem_typ = _RANDOM_848[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_fence = _RANDOM_848[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_fencei = _RANDOM_848[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_store = _RANDOM_848[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_amo = _RANDOM_848[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_load = _RANDOM_848[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_is_unique = _RANDOM_848[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_flush_on_commit = _RANDOM_848[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ldst = _RANDOM_848[19:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_lrs1 = _RANDOM_848[25:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_lrs2 = _RANDOM_848[31:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_849 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_lrs3 = _RANDOM_849[5:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_ldst_val = _RANDOM_849[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_dst_rtype = _RANDOM_849[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_lrs1_rtype = _RANDOM_849[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_lrs2_rtype = _RANDOM_849[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_frs3_en = _RANDOM_849[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_fp_val = _RANDOM_849[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_fp_single = _RANDOM_849[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_xcpt_if = _RANDOM_849[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_replay_if = _RANDOM_849[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_850 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_851 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_debug_wdata = {_RANDOM_851[17:0], _RANDOM_850, _RANDOM_849[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_852 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_18_debug_events_fetch_seq = {_RANDOM_852[17:0], _RANDOM_851[31:18]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_valid = _RANDOM_852[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_iw_state = _RANDOM_852[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_uopc = _RANDOM_852[29:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_853 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_inst = {_RANDOM_853[29:0], _RANDOM_852[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_854 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_855 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_pc = {_RANDOM_855[5:0], _RANDOM_854, _RANDOM_853[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_fu_code = _RANDOM_855[13:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_br_type = _RANDOM_855[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_op1_sel = _RANDOM_855[19:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_op2_sel = _RANDOM_855[22:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_imm_sel = _RANDOM_855[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_op_fcn = _RANDOM_855[29:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_fcn_dw = _RANDOM_855[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_rf_wen = _RANDOM_855[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_856 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_csr_cmd = _RANDOM_856[2:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_is_load = _RANDOM_856[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_is_sta = _RANDOM_856[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ctrl_is_std = _RANDOM_856[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_wakeup_delay = _RANDOM_856[7:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_allocate_brtag = _RANDOM_856[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_br_or_jmp = _RANDOM_856[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_jump = _RANDOM_856[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_jal = _RANDOM_856[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_ret = _RANDOM_856[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_call = _RANDOM_856[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_mask = _RANDOM_856[21:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_tag = _RANDOM_856[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_prediction_bpd_predict_val = _RANDOM_856[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_prediction_bpd_predict_taken = _RANDOM_856[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_prediction_btb_hit = _RANDOM_856[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_prediction_btb_predicted = _RANDOM_856[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_br_prediction_is_br_or_jalr = _RANDOM_856[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stat_brjmp_mispredicted = _RANDOM_856[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stat_btb_made_pred = _RANDOM_856[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_857 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stat_btb_mispredicted = _RANDOM_857[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stat_bpd_made_pred = _RANDOM_857[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stat_bpd_mispredicted = _RANDOM_857[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_fetch_pc_lob = _RANDOM_857[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_imm_packed = _RANDOM_857[25:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_858 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_csr_addr = {_RANDOM_858[5:0], _RANDOM_857[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_rob_idx = _RANDOM_858[11:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ldq_idx = _RANDOM_858[15:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stq_idx = _RANDOM_858[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_brob_idx = _RANDOM_858[24:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_pdst = _RANDOM_858[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_859 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_pop1 = _RANDOM_859[6:0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_pop2 = _RANDOM_859[13:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_pop3 = _RANDOM_859[20:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_prs1_busy = _RANDOM_859[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_prs2_busy = _RANDOM_859[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_prs3_busy = _RANDOM_859[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_stale_pdst = _RANDOM_859[30:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_exception = _RANDOM_859[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_860 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_861 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_exc_cause = {_RANDOM_861, _RANDOM_860};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_862 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_bypassable = _RANDOM_862[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_mem_cmd = _RANDOM_862[4:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_mem_typ = _RANDOM_862[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_fence = _RANDOM_862[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_fencei = _RANDOM_862[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_store = _RANDOM_862[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_amo = _RANDOM_862[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_load = _RANDOM_862[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_is_unique = _RANDOM_862[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_flush_on_commit = _RANDOM_862[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ldst = _RANDOM_862[20:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_lrs1 = _RANDOM_862[26:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_863 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_lrs2 = {_RANDOM_863[0], _RANDOM_862[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_lrs3 = _RANDOM_863[6:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_ldst_val = _RANDOM_863[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_dst_rtype = _RANDOM_863[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_lrs1_rtype = _RANDOM_863[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_lrs2_rtype = _RANDOM_863[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_frs3_en = _RANDOM_863[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_fp_val = _RANDOM_863[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_fp_single = _RANDOM_863[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_xcpt_if = _RANDOM_863[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_replay_if = _RANDOM_863[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_864 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_865 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_debug_wdata = {_RANDOM_865[18:0], _RANDOM_864, _RANDOM_863[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_866 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_19_debug_events_fetch_seq = {_RANDOM_866[18:0], _RANDOM_865[31:19]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_valid = _RANDOM_866[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_iw_state = _RANDOM_866[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_uopc = _RANDOM_866[30:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_867 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_inst = {_RANDOM_867[30:0], _RANDOM_866[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_868 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_869 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_pc = {_RANDOM_869[6:0], _RANDOM_868, _RANDOM_867[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_fu_code = _RANDOM_869[14:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_br_type = _RANDOM_869[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_op1_sel = _RANDOM_869[20:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_op2_sel = _RANDOM_869[23:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_imm_sel = _RANDOM_869[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_op_fcn = _RANDOM_869[30:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_fcn_dw = _RANDOM_869[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_870 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_rf_wen = _RANDOM_870[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_csr_cmd = _RANDOM_870[3:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_is_load = _RANDOM_870[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_is_sta = _RANDOM_870[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ctrl_is_std = _RANDOM_870[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_wakeup_delay = _RANDOM_870[8:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_allocate_brtag = _RANDOM_870[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_br_or_jmp = _RANDOM_870[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_jump = _RANDOM_870[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_jal = _RANDOM_870[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_ret = _RANDOM_870[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_call = _RANDOM_870[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_mask = _RANDOM_870[22:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_tag = _RANDOM_870[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_prediction_bpd_predict_val = _RANDOM_870[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_prediction_bpd_predict_taken = _RANDOM_870[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_prediction_btb_hit = _RANDOM_870[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_prediction_btb_predicted = _RANDOM_870[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_br_prediction_is_br_or_jalr = _RANDOM_870[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stat_brjmp_mispredicted = _RANDOM_870[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_871 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stat_btb_made_pred = _RANDOM_871[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stat_btb_mispredicted = _RANDOM_871[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stat_bpd_made_pred = _RANDOM_871[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stat_bpd_mispredicted = _RANDOM_871[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_fetch_pc_lob = _RANDOM_871[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_imm_packed = _RANDOM_871[26:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_872 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_csr_addr = {_RANDOM_872[6:0], _RANDOM_871[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_rob_idx = _RANDOM_872[12:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ldq_idx = _RANDOM_872[16:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stq_idx = _RANDOM_872[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_brob_idx = _RANDOM_872[25:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_873 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_pdst = {_RANDOM_873[0], _RANDOM_872[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_pop1 = _RANDOM_873[7:1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_pop2 = _RANDOM_873[14:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_pop3 = _RANDOM_873[21:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_prs1_busy = _RANDOM_873[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_prs2_busy = _RANDOM_873[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_prs3_busy = _RANDOM_873[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_stale_pdst = _RANDOM_873[31:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_874 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_exception = _RANDOM_874[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_875 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_876 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_exc_cause = {_RANDOM_876[0], _RANDOM_875, _RANDOM_874[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_bypassable = _RANDOM_876[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_mem_cmd = _RANDOM_876[5:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_mem_typ = _RANDOM_876[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_fence = _RANDOM_876[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_fencei = _RANDOM_876[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_store = _RANDOM_876[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_amo = _RANDOM_876[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_load = _RANDOM_876[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_is_unique = _RANDOM_876[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_flush_on_commit = _RANDOM_876[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ldst = _RANDOM_876[21:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_lrs1 = _RANDOM_876[27:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_877 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_lrs2 = {_RANDOM_877[1:0], _RANDOM_876[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_lrs3 = _RANDOM_877[7:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_ldst_val = _RANDOM_877[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_dst_rtype = _RANDOM_877[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_lrs1_rtype = _RANDOM_877[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_lrs2_rtype = _RANDOM_877[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_frs3_en = _RANDOM_877[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_fp_val = _RANDOM_877[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_fp_single = _RANDOM_877[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_xcpt_if = _RANDOM_877[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_replay_if = _RANDOM_877[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_878 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_879 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_debug_wdata = {_RANDOM_879[19:0], _RANDOM_878, _RANDOM_877[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_880 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_20_debug_events_fetch_seq = {_RANDOM_880[19:0], _RANDOM_879[31:20]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_valid = _RANDOM_880[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_iw_state = _RANDOM_880[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_uopc = _RANDOM_880[31:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_881 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_inst = _RANDOM_881;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_882 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_883 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_pc = {_RANDOM_883[7:0], _RANDOM_882};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_fu_code = _RANDOM_883[15:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_br_type = _RANDOM_883[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_op1_sel = _RANDOM_883[21:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_op2_sel = _RANDOM_883[24:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_imm_sel = _RANDOM_883[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_op_fcn = _RANDOM_883[31:28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_884 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_fcn_dw = _RANDOM_884[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_rf_wen = _RANDOM_884[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_csr_cmd = _RANDOM_884[4:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_is_load = _RANDOM_884[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_is_sta = _RANDOM_884[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ctrl_is_std = _RANDOM_884[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_wakeup_delay = _RANDOM_884[9:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_allocate_brtag = _RANDOM_884[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_br_or_jmp = _RANDOM_884[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_jump = _RANDOM_884[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_jal = _RANDOM_884[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_ret = _RANDOM_884[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_call = _RANDOM_884[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_mask = _RANDOM_884[23:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_tag = _RANDOM_884[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_prediction_bpd_predict_val = _RANDOM_884[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_prediction_bpd_predict_taken = _RANDOM_884[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_prediction_btb_hit = _RANDOM_884[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_prediction_btb_predicted = _RANDOM_884[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_br_prediction_is_br_or_jalr = _RANDOM_884[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_885 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stat_brjmp_mispredicted = _RANDOM_885[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stat_btb_made_pred = _RANDOM_885[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stat_btb_mispredicted = _RANDOM_885[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stat_bpd_made_pred = _RANDOM_885[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stat_bpd_mispredicted = _RANDOM_885[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_fetch_pc_lob = _RANDOM_885[7:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_imm_packed = _RANDOM_885[27:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_886 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_csr_addr = {_RANDOM_886[7:0], _RANDOM_885[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_rob_idx = _RANDOM_886[13:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ldq_idx = _RANDOM_886[17:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stq_idx = _RANDOM_886[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_brob_idx = _RANDOM_886[26:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_887 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_pdst = {_RANDOM_887[1:0], _RANDOM_886[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_pop1 = _RANDOM_887[8:2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_pop2 = _RANDOM_887[15:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_pop3 = _RANDOM_887[22:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_prs1_busy = _RANDOM_887[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_prs2_busy = _RANDOM_887[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_prs3_busy = _RANDOM_887[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_888 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_stale_pdst = {_RANDOM_888[0], _RANDOM_887[31:26]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_exception = _RANDOM_888[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_889 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_890 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_exc_cause = {_RANDOM_890[1:0], _RANDOM_889, _RANDOM_888[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_bypassable = _RANDOM_890[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_mem_cmd = _RANDOM_890[6:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_mem_typ = _RANDOM_890[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_fence = _RANDOM_890[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_fencei = _RANDOM_890[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_store = _RANDOM_890[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_amo = _RANDOM_890[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_load = _RANDOM_890[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_is_unique = _RANDOM_890[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_flush_on_commit = _RANDOM_890[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ldst = _RANDOM_890[22:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_lrs1 = _RANDOM_890[28:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_891 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_lrs2 = {_RANDOM_891[2:0], _RANDOM_890[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_lrs3 = _RANDOM_891[8:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_ldst_val = _RANDOM_891[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_dst_rtype = _RANDOM_891[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_lrs1_rtype = _RANDOM_891[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_lrs2_rtype = _RANDOM_891[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_frs3_en = _RANDOM_891[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_fp_val = _RANDOM_891[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_fp_single = _RANDOM_891[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_xcpt_if = _RANDOM_891[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_replay_if = _RANDOM_891[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_892 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_893 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_debug_wdata = {_RANDOM_893[20:0], _RANDOM_892, _RANDOM_891[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_894 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_21_debug_events_fetch_seq = {_RANDOM_894[20:0], _RANDOM_893[31:21]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_valid = _RANDOM_894[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_iw_state = _RANDOM_894[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_895 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_uopc = {_RANDOM_895[0], _RANDOM_894[31:24]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_896 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_inst = {_RANDOM_896[0], _RANDOM_895[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_897 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_pc = {_RANDOM_897[8:0], _RANDOM_896[31:1]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_fu_code = _RANDOM_897[16:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_br_type = _RANDOM_897[20:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_op1_sel = _RANDOM_897[22:21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_op2_sel = _RANDOM_897[25:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_imm_sel = _RANDOM_897[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_898 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_op_fcn = {_RANDOM_898[0], _RANDOM_897[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_fcn_dw = _RANDOM_898[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_rf_wen = _RANDOM_898[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_csr_cmd = _RANDOM_898[5:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_is_load = _RANDOM_898[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_is_sta = _RANDOM_898[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ctrl_is_std = _RANDOM_898[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_wakeup_delay = _RANDOM_898[10:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_allocate_brtag = _RANDOM_898[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_br_or_jmp = _RANDOM_898[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_jump = _RANDOM_898[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_jal = _RANDOM_898[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_ret = _RANDOM_898[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_call = _RANDOM_898[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_mask = _RANDOM_898[24:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_tag = _RANDOM_898[27:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_prediction_bpd_predict_val = _RANDOM_898[28];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_prediction_bpd_predict_taken = _RANDOM_898[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_prediction_btb_hit = _RANDOM_898[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_prediction_btb_predicted = _RANDOM_898[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_899 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_br_prediction_is_br_or_jalr = _RANDOM_899[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stat_brjmp_mispredicted = _RANDOM_899[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stat_btb_made_pred = _RANDOM_899[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stat_btb_mispredicted = _RANDOM_899[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stat_bpd_made_pred = _RANDOM_899[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stat_bpd_mispredicted = _RANDOM_899[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_fetch_pc_lob = _RANDOM_899[8:6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_imm_packed = _RANDOM_899[28:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_900 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_csr_addr = {_RANDOM_900[8:0], _RANDOM_899[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_rob_idx = _RANDOM_900[14:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ldq_idx = _RANDOM_900[18:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stq_idx = _RANDOM_900[22:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_brob_idx = _RANDOM_900[27:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_901 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_pdst = {_RANDOM_901[2:0], _RANDOM_900[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_pop1 = _RANDOM_901[9:3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_pop2 = _RANDOM_901[16:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_pop3 = _RANDOM_901[23:17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_prs1_busy = _RANDOM_901[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_prs2_busy = _RANDOM_901[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_prs3_busy = _RANDOM_901[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_902 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_stale_pdst = {_RANDOM_902[1:0], _RANDOM_901[31:27]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_exception = _RANDOM_902[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_903 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_904 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_exc_cause = {_RANDOM_904[2:0], _RANDOM_903, _RANDOM_902[31:3]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_bypassable = _RANDOM_904[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_mem_cmd = _RANDOM_904[7:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_mem_typ = _RANDOM_904[10:8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_fence = _RANDOM_904[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_fencei = _RANDOM_904[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_store = _RANDOM_904[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_amo = _RANDOM_904[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_load = _RANDOM_904[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_is_unique = _RANDOM_904[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_flush_on_commit = _RANDOM_904[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ldst = _RANDOM_904[23:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_lrs1 = _RANDOM_904[29:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_905 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_lrs2 = {_RANDOM_905[3:0], _RANDOM_904[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_lrs3 = _RANDOM_905[9:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_ldst_val = _RANDOM_905[10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_dst_rtype = _RANDOM_905[12:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_lrs1_rtype = _RANDOM_905[14:13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_lrs2_rtype = _RANDOM_905[16:15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_frs3_en = _RANDOM_905[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_fp_val = _RANDOM_905[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_fp_single = _RANDOM_905[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_xcpt_if = _RANDOM_905[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_replay_if = _RANDOM_905[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_906 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_907 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_debug_wdata = {_RANDOM_907[21:0], _RANDOM_906, _RANDOM_905[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_908 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_22_debug_events_fetch_seq = {_RANDOM_908[21:0], _RANDOM_907[31:22]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_valid = _RANDOM_908[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_iw_state = _RANDOM_908[24:23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_909 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_uopc = {_RANDOM_909[1:0], _RANDOM_908[31:25]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_910 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_inst = {_RANDOM_910[1:0], _RANDOM_909[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_911 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_pc = {_RANDOM_911[9:0], _RANDOM_910[31:2]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_fu_code = _RANDOM_911[17:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_br_type = _RANDOM_911[21:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_op1_sel = _RANDOM_911[23:22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_op2_sel = _RANDOM_911[26:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_imm_sel = _RANDOM_911[29:27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_912 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_op_fcn = {_RANDOM_912[1:0], _RANDOM_911[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_fcn_dw = _RANDOM_912[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_rf_wen = _RANDOM_912[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_csr_cmd = _RANDOM_912[6:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_is_load = _RANDOM_912[7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_is_sta = _RANDOM_912[8];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ctrl_is_std = _RANDOM_912[9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_wakeup_delay = _RANDOM_912[11:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_allocate_brtag = _RANDOM_912[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_br_or_jmp = _RANDOM_912[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_jump = _RANDOM_912[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_jal = _RANDOM_912[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_ret = _RANDOM_912[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_call = _RANDOM_912[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_mask = _RANDOM_912[25:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_tag = _RANDOM_912[28:26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_prediction_bpd_predict_val = _RANDOM_912[29];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_prediction_bpd_predict_taken = _RANDOM_912[30];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_prediction_btb_hit = _RANDOM_912[31];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_913 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_prediction_btb_predicted = _RANDOM_913[0];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_br_prediction_is_br_or_jalr = _RANDOM_913[1];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stat_brjmp_mispredicted = _RANDOM_913[2];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stat_btb_made_pred = _RANDOM_913[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stat_btb_mispredicted = _RANDOM_913[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stat_bpd_made_pred = _RANDOM_913[5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stat_bpd_mispredicted = _RANDOM_913[6];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_fetch_pc_lob = _RANDOM_913[9:7];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_imm_packed = _RANDOM_913[29:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_914 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_csr_addr = {_RANDOM_914[9:0], _RANDOM_913[31:30]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_rob_idx = _RANDOM_914[15:10];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ldq_idx = _RANDOM_914[19:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stq_idx = _RANDOM_914[23:20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_brob_idx = _RANDOM_914[28:24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_915 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_pdst = {_RANDOM_915[3:0], _RANDOM_914[31:29]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_pop1 = _RANDOM_915[10:4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_pop2 = _RANDOM_915[17:11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_pop3 = _RANDOM_915[24:18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_prs1_busy = _RANDOM_915[25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_prs2_busy = _RANDOM_915[26];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_prs3_busy = _RANDOM_915[27];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_916 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_stale_pdst = {_RANDOM_916[2:0], _RANDOM_915[31:28]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_exception = _RANDOM_916[3];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_917 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_918 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_exc_cause = {_RANDOM_918[3:0], _RANDOM_917, _RANDOM_916[31:4]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_bypassable = _RANDOM_918[4];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_mem_cmd = _RANDOM_918[8:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_mem_typ = _RANDOM_918[11:9];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_fence = _RANDOM_918[12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_fencei = _RANDOM_918[13];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_store = _RANDOM_918[14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_amo = _RANDOM_918[15];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_load = _RANDOM_918[16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_is_unique = _RANDOM_918[17];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_flush_on_commit = _RANDOM_918[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ldst = _RANDOM_918[24:19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_lrs1 = _RANDOM_918[30:25];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_919 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_lrs2 = {_RANDOM_919[4:0], _RANDOM_918[31]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_lrs3 = _RANDOM_919[10:5];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_ldst_val = _RANDOM_919[11];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_dst_rtype = _RANDOM_919[13:12];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_lrs1_rtype = _RANDOM_919[15:14];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_lrs2_rtype = _RANDOM_919[17:16];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_frs3_en = _RANDOM_919[18];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_fp_val = _RANDOM_919[19];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_fp_single = _RANDOM_919[20];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_xcpt_if = _RANDOM_919[21];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_replay_if = _RANDOM_919[22];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_920 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_921 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_debug_wdata = {_RANDOM_921[22:0], _RANDOM_920, _RANDOM_919[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        _RANDOM_922 = `RANDOM;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_38110_23_debug_events_fetch_seq = {_RANDOM_922[22:0], _RANDOM_921[31:23]};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1557:5
        T_47576 = _RANDOM_922[23];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2940:5
        T_47616 = _RANDOM_922[24];	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2978:5
      `endif
    end // initial
  `endif
      wire _T_47631 = _T_3 & casez_tmp_76;	// rob.scala:453:59, :624:41
      wire _T_47632 = casez_tmp_64 | casez_tmp_62;	// rob.scala:453:59, :626:48
      wire _T_47635 = _T_47631 & ~_T_47632;	// rob.scala:625:46, :626:23
      wire _T_47660 = _T_4 & casez_tmp_168;	// rob.scala:453:59, :624:41
      wire _T_47661 = casez_tmp_156 | casez_tmp_154;	// rob.scala:453:59, :626:48
      wire _T_47664 = _T_47660 & ~_T_47661;	// rob.scala:625:46, :626:23
      wire [1:0] _T_48125 = {casez_tmp_94, casez_tmp_2};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:3152:20, rob.scala:433:51
      wire _T_48130 = rob_head == rob_tail;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :717:59
  assign _T = |{_T_4, _T_3} & ({_T_4, _T_3} ^ _T_48125) == 2'h0 & ~(r_partial_row & _T_48130);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:59, :3149:20, :3151:20, rob.scala:301:21, :715:53, :716:{52,76,89}, :717:{31,47}
      wire _T_48185 = rob_tail == 5'h17;	// rob.scala:192:32, :347:34, util.scala:75:28
      wire _T_48195 = _T_48130 & _T_48125 == 2'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:59, rob.scala:759:{40,65}
      wire [63:0] _T_6 = {24'h0, r_xcpt_badvaddr};	// Bitwise.scala:33:12, rob.scala:882:27, util.scala:114:43
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_0_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_185 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_185 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_185 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_185 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_0_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_186 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_186 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_186 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_186 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_1_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_187 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_187 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_187 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_187 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_1_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_188 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_188 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_188 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_188 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_2_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_189 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_189 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_189 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_189 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_2_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_190 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_190 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_190 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_190 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_3_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_191 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_191 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_191 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_191 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_3_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_192 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_192 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_192 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_192 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_4_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_193 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_193 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_193 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_193 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_4_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_194 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_194 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_194 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_194 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_5_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_195 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_195 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_195 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_195 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_5_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_196 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_196 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_196 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_196 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_6_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_197 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_197 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_197 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_197 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_6_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_198 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_198 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_198 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_198 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_7_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_199 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_199 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_199 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_199 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_7_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_200 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_200 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_200 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_200 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_8_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_201 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_201 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_201 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_201 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_8_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_202 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_202 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_202 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_202 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_9_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_203 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_203 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_203 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_203 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_9_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_204 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_204 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_204 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_204 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_10_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_205 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_205 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_205 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_205 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_10_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_206 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_206 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_206 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_206 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_11_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_207 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_207 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_207 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_207 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_11_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_208 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_208 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_208 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_208 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_12_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_209 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_209 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_209 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_209 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_12_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_210 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_210 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_210 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_210 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_13_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_211 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_211 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_211 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_211 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_13_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_212 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_212 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_212 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_212 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_14_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_213 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_213 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_213 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_213 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_14_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_214 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_214 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_214 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_214 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_15_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_215 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_215 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_215 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_215 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_15_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_216 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_216 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_216 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_216 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_16_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_217 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_217 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_217 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_217 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_16_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_218 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_218 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_218 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_218 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_17_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_219 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_219 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_219 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_219 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_17_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_220 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_220 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_220 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_220 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_18_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_221 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_221 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_221 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_221 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_18_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_222 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_222 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_222 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_222 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_19_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_223 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_223 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_223 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_223 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_19_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_224 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_224 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_224 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_224 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_20_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_225 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_225 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_225 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_225 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_20_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_226 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_226 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_226 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_226 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_21_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_227 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_227 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_227 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_227 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_21_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_228 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_228 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_228 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_228 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_22_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_229 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_229 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_229 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_229 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_22_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_230 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_230 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_230 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_230 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_26182_23_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_231 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_231 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_231 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_231 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
  always @(*) begin	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    casez (T_38110_23_dst_rtype)	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b00:
        casez_tmp_232 = 8'h58;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b01:
        casez_tmp_232 = 8'h66;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      2'b10:
        casez_tmp_232 = 8'h2D;	// rob.scala:946:18, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
      default:
        casez_tmp_232 = 8'h43;	// rob.scala:1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
    endcase	// rob.scala:350:34, :1048:{21,58}, :1049:{21,58}, :1050:{21,58}, :1051:{21,58}
  end // always @(*)
      wire _T_48144 = _T_29097 & rob_tail != rob_head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :726:{35,47}
      wire [1:0] _T_7 = rob_state == 2'h0 ? 2'h1 : rob_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:59, Conditional.scala:24:42, rob.scala:443:23, :453:100, :777:23
      wire [1:0] _T_8 = rob_state == 2'h2 & _T_48195 ? 2'h1 : rob_state == 2'h1 ? (_T_47568 ? 2'h2 : _T_23671 |
                _T_23670 ? 2'h3 : _T_47568 ? 2'h2 : _T_7) : _T_7;	// Conditional.scala:24:42, rob.scala:443:23, :453:100, :783:26, :791:32, :800:26, :931:42
      wire _T_32357 = ~(io_wb_resps_0_valid & ~_T_28590 & ~casez_tmp_84) | reset;	// rob.scala:331:55, :535:{17,18,75}, :536:22
      wire _T_32369 = ~(io_wb_resps_0_valid & ~_T_28590 & casez_tmp_86 & casez_tmp_85 !=
                io_wb_resps_0_bits_uop_pdst) | reset;	// rob.scala:331:55, :538:{17,18,75}, :539:{37,54}
      wire _T_32561 = ~(io_wb_resps_1_valid & ~_T_28598 & ~casez_tmp_87) | reset;	// rob.scala:331:55, :535:{17,18,75}, :536:22
      wire _T_32573 = ~(io_wb_resps_1_valid & ~_T_28598 & casez_tmp_89 & casez_tmp_88 !=
                io_wb_resps_1_bits_uop_pdst) | reset;	// rob.scala:331:55, :538:{17,18,75}, :539:{37,54}
      wire _T_32765 = ~(io_wb_resps_2_valid & ~_T_28606 & ~casez_tmp_90) | reset;	// rob.scala:331:55, :535:{17,18,75}, :536:22
      wire _T_32777 = ~(io_wb_resps_2_valid & ~_T_28606 & casez_tmp_92 & casez_tmp_91 !=
                io_wb_resps_2_bits_uop_pdst) | reset;	// rob.scala:331:55, :538:{17,18,75}, :539:{37,54}
      wire _T_44285 = ~(io_wb_resps_0_valid & _T_28590 & ~casez_tmp_176) | reset;	// rob.scala:535:{17,18,75}, :536:22
      wire _T_44297 = ~(io_wb_resps_0_valid & _T_28590 & casez_tmp_178 & casez_tmp_177 !=
                io_wb_resps_0_bits_uop_pdst) | reset;	// rob.scala:538:{17,18,75}, :539:{37,54}
      wire _T_44489 = ~(io_wb_resps_1_valid & _T_28598 & ~casez_tmp_179) | reset;	// rob.scala:535:{17,18,75}, :536:22
      wire _T_44501 = ~(io_wb_resps_1_valid & _T_28598 & casez_tmp_181 & casez_tmp_180 !=
                io_wb_resps_1_bits_uop_pdst) | reset;	// rob.scala:538:{17,18,75}, :539:{37,54}
      wire _T_44693 = ~(io_wb_resps_2_valid & _T_28606 & ~casez_tmp_182) | reset;	// rob.scala:535:{17,18,75}, :536:22
      wire _T_44705 = ~(io_wb_resps_2_valid & _T_28606 & casez_tmp_184 & casez_tmp_183 !=
                io_wb_resps_2_bits_uop_pdst) | reset;	// rob.scala:538:{17,18,75}, :539:{37,54}
      wire _T_47646 = ~(_T_3 & ~casez_tmp_76 & |T_28314_R0_data) | reset;	// rob.scala:340:30, :453:59, :630:{14,15}, :631:{16,39}, :632:35
      wire _T_47657 = ~(_T_47631 & _T_47632 & |T_28314_R0_data) | reset;	// rob.scala:340:30, :632:35, :634:{14,15}, :636:68
      wire _T_47675 = ~(_T_4 & ~casez_tmp_168 & |T_40242_R0_data) | reset;	// rob.scala:340:30, :453:59, :630:{14,15}, :631:{16,39}, :632:35
      wire _T_47686 = ~(_T_47660 & _T_47661 & |T_40242_R0_data) | reset;	// rob.scala:340:30, :632:35, :634:{14,15}, :636:68
      wire _T_48314 = rob_head == 5'h1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48316 = rob_tail == 5'h1;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48400 = rob_head == 5'h2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48402 = rob_tail == 5'h2;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48486 = rob_head == 5'h3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48488 = rob_tail == 5'h3;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48572 = rob_head == 5'h4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48574 = rob_tail == 5'h4;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48658 = rob_head == 5'h5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48660 = rob_tail == 5'h5;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48744 = rob_head == 5'h6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48746 = rob_tail == 5'h6;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48830 = rob_head == 5'h7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48832 = rob_tail == 5'h7;	// rob.scala:192:32, :347:34, :970:50
      wire _T_48916 = rob_head == 5'h8;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48918 = rob_tail == 5'h8;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49002 = rob_head == 5'h9;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49004 = rob_tail == 5'h9;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49088 = rob_head == 5'hA;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49090 = rob_tail == 5'hA;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49174 = rob_head == 5'hB;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49176 = rob_tail == 5'hB;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49260 = rob_head == 5'hC;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49262 = rob_tail == 5'hC;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49346 = rob_head == 5'hD;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49348 = rob_tail == 5'hD;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49432 = rob_head == 5'hE;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49434 = rob_tail == 5'hE;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49518 = rob_head == 5'hF;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49520 = rob_tail == 5'hF;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49604 = rob_head == 5'h10;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49606 = rob_tail == 5'h10;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49690 = rob_head == 5'h11;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49692 = rob_tail == 5'h11;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49776 = rob_head == 5'h12;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49778 = rob_tail == 5'h12;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49862 = rob_head == 5'h13;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49864 = rob_tail == 5'h13;	// rob.scala:192:32, :347:34, :970:50
      wire _T_49948 = rob_head == 5'h14;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_49950 = rob_tail == 5'h14;	// rob.scala:192:32, :347:34, :970:50
      wire _T_50034 = rob_head == 5'h15;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_50036 = rob_tail == 5'h15;	// rob.scala:192:32, :347:34, :970:50
      wire _T_50120 = rob_head == 5'h16;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_50122 = rob_tail == 5'h16;	// rob.scala:192:32, :347:34, :970:50
      wire _T_50206 = rob_head == 5'h17;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :970:26
      wire _T_48103 = ~(_T_47568 & ~io_cxcpt_valid & ~r_xcpt_val) | reset;	// rob.scala:667:16, :693:{11,12,34,50,53}
      wire _T_48109 = ~(_T_48195 & r_xcpt_val) | reset;	// rob.scala:667:16, :696:{11,12,23}
      wire _T_48118 = ~(_will_throw_exception & r_xcpt_uop_rob_idx[5:1] != rob_head) | reset;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:222:27, :650:80, :699:{11,12,35,69}
      wire [5:0] _rob_tail_idx = {rob_tail, 1'h0};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:192:32
      wire _T_9 = rob_tail == 5'h1;	// rob.scala:192:32, :347:34
      wire _T_10 = rob_tail == 5'h2;	// rob.scala:192:32, :347:34
      wire _T_11 = rob_tail == 5'h3;	// rob.scala:192:32, :347:34
      wire _T_12 = rob_tail == 5'h4;	// rob.scala:192:32, :347:34
      wire _T_13 = rob_tail == 5'h5;	// rob.scala:192:32, :347:34
      wire _T_14 = rob_tail == 5'h6;	// rob.scala:192:32, :347:34
      wire _T_15 = rob_tail == 5'h7;	// rob.scala:192:32, :347:34
      wire _T_16 = rob_tail == 5'h8;	// rob.scala:192:32, :347:34
      wire _T_17 = rob_tail == 5'h9;	// rob.scala:192:32, :347:34
      wire _T_18 = rob_tail == 5'hA;	// rob.scala:192:32, :347:34
      wire _T_19 = rob_tail == 5'hB;	// rob.scala:192:32, :347:34
      wire _T_20 = rob_tail == 5'hC;	// rob.scala:192:32, :347:34
      wire _T_21 = rob_tail == 5'hD;	// rob.scala:192:32, :347:34
      wire _T_22 = rob_tail == 5'hE;	// rob.scala:192:32, :347:34
      wire _T_23 = rob_tail == 5'hF;	// rob.scala:192:32, :347:34
      wire _T_24 = rob_tail == 5'h10;	// rob.scala:192:32, :347:34
      wire _T_25 = rob_tail == 5'h11;	// rob.scala:192:32, :347:34
      wire _T_26 = rob_tail == 5'h12;	// rob.scala:192:32, :347:34
      wire _T_27 = rob_tail == 5'h13;	// rob.scala:192:32, :347:34
      wire _T_28 = rob_tail == 5'h14;	// rob.scala:192:32, :347:34
      wire _T_29 = rob_tail == 5'h15;	// rob.scala:192:32, :347:34
      wire _T_30 = rob_tail == 5'h16;	// rob.scala:192:32, :347:34
      wire _T_31 = rob_tail == 5'h17;	// rob.scala:192:32, :347:34
      wire [31:0] _T_32 = ~io_dis_valids_0 | |rob_tail ? T_26182_0_inst : io_dis_uops_0_inst;	// rob.scala:192:32, :347:34, :350:34
      wire [31:0] _T_33 = io_dis_valids_0 & _T_9 ? io_dis_uops_0_inst : T_26182_1_inst;	// rob.scala:350:34
      wire [31:0] _T_34 = io_dis_valids_0 & _T_10 ? io_dis_uops_0_inst : T_26182_2_inst;	// rob.scala:350:34
      wire [31:0] _T_35 = io_dis_valids_0 & _T_11 ? io_dis_uops_0_inst : T_26182_3_inst;	// rob.scala:350:34
      wire [31:0] _T_36 = io_dis_valids_0 & _T_12 ? io_dis_uops_0_inst : T_26182_4_inst;	// rob.scala:350:34
      wire [31:0] _T_37 = io_dis_valids_0 & _T_13 ? io_dis_uops_0_inst : T_26182_5_inst;	// rob.scala:350:34
      wire [31:0] _T_38 = io_dis_valids_0 & _T_14 ? io_dis_uops_0_inst : T_26182_6_inst;	// rob.scala:350:34
      wire [31:0] _T_39 = io_dis_valids_0 & _T_15 ? io_dis_uops_0_inst : T_26182_7_inst;	// rob.scala:350:34
      wire [31:0] _T_40 = io_dis_valids_0 & _T_16 ? io_dis_uops_0_inst : T_26182_8_inst;	// rob.scala:350:34
      wire [31:0] _T_41 = io_dis_valids_0 & _T_17 ? io_dis_uops_0_inst : T_26182_9_inst;	// rob.scala:350:34
      wire [31:0] _T_42 = io_dis_valids_0 & _T_18 ? io_dis_uops_0_inst : T_26182_10_inst;	// rob.scala:350:34
      wire [31:0] _T_43 = io_dis_valids_0 & _T_19 ? io_dis_uops_0_inst : T_26182_11_inst;	// rob.scala:350:34
      wire [31:0] _T_44 = io_dis_valids_0 & _T_20 ? io_dis_uops_0_inst : T_26182_12_inst;	// rob.scala:350:34
      wire [31:0] _T_45 = io_dis_valids_0 & _T_21 ? io_dis_uops_0_inst : T_26182_13_inst;	// rob.scala:350:34
      wire [31:0] _T_46 = io_dis_valids_0 & _T_22 ? io_dis_uops_0_inst : T_26182_14_inst;	// rob.scala:350:34
      wire [31:0] _T_47 = io_dis_valids_0 & _T_23 ? io_dis_uops_0_inst : T_26182_15_inst;	// rob.scala:350:34
      wire [31:0] _T_48 = io_dis_valids_0 & _T_24 ? io_dis_uops_0_inst : T_26182_16_inst;	// rob.scala:350:34
      wire [31:0] _T_49 = io_dis_valids_0 & _T_25 ? io_dis_uops_0_inst : T_26182_17_inst;	// rob.scala:350:34
      wire [31:0] _T_50 = io_dis_valids_0 & _T_26 ? io_dis_uops_0_inst : T_26182_18_inst;	// rob.scala:350:34
      wire [31:0] _T_51 = io_dis_valids_0 & _T_27 ? io_dis_uops_0_inst : T_26182_19_inst;	// rob.scala:350:34
      wire [31:0] _T_52 = io_dis_valids_0 & _T_28 ? io_dis_uops_0_inst : T_26182_20_inst;	// rob.scala:350:34
      wire [31:0] _T_53 = io_dis_valids_0 & _T_29 ? io_dis_uops_0_inst : T_26182_21_inst;	// rob.scala:350:34
      wire [31:0] _T_54 = io_dis_valids_0 & _T_30 ? io_dis_uops_0_inst : T_26182_22_inst;	// rob.scala:350:34
      wire [31:0] _T_55 = io_dis_valids_0 & _T_31 ? io_dis_uops_0_inst : T_26182_23_inst;	// rob.scala:350:34
      wire _T_56 = ~io_dis_valids_0 & _T_23559 & ~casez_tmp;	// rob.scala:346:7, :355:47, :356:7
      wire _T_28620 = io_brinfo_rob_idx[0];	// rob.scala:227:38
      wire _T_28623 = io_brinfo_valid & ~_T_28620;	// rob.scala:331:55, :400:29
      wire [4:0] _io_brinfo_rob_idx_5to1 = io_brinfo_rob_idx[5:1];	// rob.scala:222:27
      wire _T_57 = _io_brinfo_rob_idx_5to1 == 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, rob.scala:402:72
      wire _T_58 = _io_brinfo_rob_idx_5to1 == 5'h1;	// rob.scala:347:34, :402:72
      wire _T_59 = _io_brinfo_rob_idx_5to1 == 5'h2;	// rob.scala:347:34, :402:72
      wire _T_60 = _io_brinfo_rob_idx_5to1 == 5'h3;	// rob.scala:347:34, :402:72
      wire _T_61 = _io_brinfo_rob_idx_5to1 == 5'h4;	// rob.scala:347:34, :402:72
      wire _T_62 = _io_brinfo_rob_idx_5to1 == 5'h5;	// rob.scala:347:34, :402:72
      wire _T_63 = _io_brinfo_rob_idx_5to1 == 5'h6;	// rob.scala:347:34, :402:72
      wire _T_64 = _io_brinfo_rob_idx_5to1 == 5'h7;	// rob.scala:347:34, :402:72
      wire _T_65 = _io_brinfo_rob_idx_5to1 == 5'h8;	// rob.scala:347:34, :402:72
      wire _T_66 = _io_brinfo_rob_idx_5to1 == 5'h9;	// rob.scala:347:34, :402:72
      wire _T_67 = _io_brinfo_rob_idx_5to1 == 5'hA;	// rob.scala:347:34, :402:72
      wire _T_68 = _io_brinfo_rob_idx_5to1 == 5'hB;	// rob.scala:347:34, :402:72
      wire _T_69 = _io_brinfo_rob_idx_5to1 == 5'hC;	// rob.scala:347:34, :402:72
      wire _T_70 = _io_brinfo_rob_idx_5to1 == 5'hD;	// rob.scala:347:34, :402:72
      wire _T_71 = _io_brinfo_rob_idx_5to1 == 5'hE;	// rob.scala:347:34, :402:72
      wire _T_72 = _io_brinfo_rob_idx_5to1 == 5'hF;	// rob.scala:347:34, :402:72
      wire _T_73 = _io_brinfo_rob_idx_5to1 == 5'h10;	// rob.scala:347:34, :402:72
      wire _T_74 = _io_brinfo_rob_idx_5to1 == 5'h11;	// rob.scala:347:34, :402:72
      wire _T_75 = _io_brinfo_rob_idx_5to1 == 5'h12;	// rob.scala:347:34, :402:72
      wire _T_76 = _io_brinfo_rob_idx_5to1 == 5'h13;	// rob.scala:347:34, :402:72
      wire _T_77 = _io_brinfo_rob_idx_5to1 == 5'h14;	// rob.scala:347:34, :402:72
      wire _T_78 = _io_brinfo_rob_idx_5to1 == 5'h15;	// rob.scala:347:34, :402:72
      wire _T_79 = _io_brinfo_rob_idx_5to1 == 5'h16;	// rob.scala:347:34, :402:72
      wire _T_80 = _io_brinfo_rob_idx_5to1 == 5'h17;	// rob.scala:347:34, :402:72
      wire _T_81 = rob_head == 5'h1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_82 = rob_head == 5'h2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_83 = rob_head == 5'h3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_84 = rob_head == 5'h4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_85 = rob_head == 5'h5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_86 = rob_head == 5'h6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_87 = rob_head == 5'h7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_88 = rob_head == 5'h8;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_89 = rob_head == 5'h9;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_90 = rob_head == 5'hA;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_91 = rob_head == 5'hB;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_92 = rob_head == 5'hC;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_93 = rob_head == 5'hD;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_94 = rob_head == 5'hE;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_95 = rob_head == 5'hF;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_96 = rob_head == 5'h10;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_97 = rob_head == 5'h11;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_98 = rob_head == 5'h12;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_99 = rob_head == 5'h13;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_100 = rob_head == 5'h14;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_101 = rob_head == 5'h15;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_102 = rob_head == 5'h16;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_103 = rob_head == 5'h17;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:347:34, :433:51
      wire _T_29368 = T_23706_0 & |(io_brinfo_mask & T_26182_0_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29369 = io_brinfo_valid & io_brinfo_mispredict;	// rob.scala:484:32
      wire _T_29370 = _T_29369 & _T_29368;	// rob.scala:484:56
      wire _T_104 = _T_29370 | ~(~_T_56 | |rob_tail);	// rob.scala:192:32, :347:34, :357:33, :487:35
      wire _T_29470 = T_23706_1 & |(io_brinfo_mask & T_26182_1_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29472 = _T_29369 & _T_29470;	// rob.scala:484:56
      wire _T_105 = _T_29472 | _T_56 & _T_9;	// rob.scala:357:33, :487:35
      wire _T_29572 = T_23706_2 & |(io_brinfo_mask & T_26182_2_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29574 = _T_29369 & _T_29572;	// rob.scala:484:56
      wire _T_106 = _T_29574 | _T_56 & _T_10;	// rob.scala:357:33, :487:35
      wire _T_29674 = T_23706_3 & |(io_brinfo_mask & T_26182_3_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29676 = _T_29369 & _T_29674;	// rob.scala:484:56
      wire _T_107 = _T_29676 | _T_56 & _T_11;	// rob.scala:357:33, :487:35
      wire _T_29776 = T_23706_4 & |(io_brinfo_mask & T_26182_4_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29778 = _T_29369 & _T_29776;	// rob.scala:484:56
      wire _T_108 = _T_29778 | _T_56 & _T_12;	// rob.scala:357:33, :487:35
      wire _T_29878 = T_23706_5 & |(io_brinfo_mask & T_26182_5_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29880 = _T_29369 & _T_29878;	// rob.scala:484:56
      wire _T_109 = _T_29880 | _T_56 & _T_13;	// rob.scala:357:33, :487:35
      wire _T_29980 = T_23706_6 & |(io_brinfo_mask & T_26182_6_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_29982 = _T_29369 & _T_29980;	// rob.scala:484:56
      wire _T_110 = _T_29982 | _T_56 & _T_14;	// rob.scala:357:33, :487:35
      wire _T_30082 = T_23706_7 & |(io_brinfo_mask & T_26182_7_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30084 = _T_29369 & _T_30082;	// rob.scala:484:56
      wire _T_111 = _T_30084 | _T_56 & _T_15;	// rob.scala:357:33, :487:35
      wire _T_30184 = T_23706_8 & |(io_brinfo_mask & T_26182_8_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30186 = _T_29369 & _T_30184;	// rob.scala:484:56
      wire _T_112 = _T_30186 | _T_56 & _T_16;	// rob.scala:357:33, :487:35
      wire _T_30286 = T_23706_9 & |(io_brinfo_mask & T_26182_9_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30288 = _T_29369 & _T_30286;	// rob.scala:484:56
      wire _T_113 = _T_30288 | _T_56 & _T_17;	// rob.scala:357:33, :487:35
      wire _T_30388 = T_23706_10 & |(io_brinfo_mask & T_26182_10_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30390 = _T_29369 & _T_30388;	// rob.scala:484:56
      wire _T_114 = _T_30390 | _T_56 & _T_18;	// rob.scala:357:33, :487:35
      wire _T_30490 = T_23706_11 & |(io_brinfo_mask & T_26182_11_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30492 = _T_29369 & _T_30490;	// rob.scala:484:56
      wire _T_115 = _T_30492 | _T_56 & _T_19;	// rob.scala:357:33, :487:35
      wire _T_30592 = T_23706_12 & |(io_brinfo_mask & T_26182_12_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30594 = _T_29369 & _T_30592;	// rob.scala:484:56
      wire _T_116 = _T_30594 | _T_56 & _T_20;	// rob.scala:357:33, :487:35
      wire _T_30694 = T_23706_13 & |(io_brinfo_mask & T_26182_13_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30696 = _T_29369 & _T_30694;	// rob.scala:484:56
      wire _T_117 = _T_30696 | _T_56 & _T_21;	// rob.scala:357:33, :487:35
      wire _T_30796 = T_23706_14 & |(io_brinfo_mask & T_26182_14_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30798 = _T_29369 & _T_30796;	// rob.scala:484:56
      wire _T_118 = _T_30798 | _T_56 & _T_22;	// rob.scala:357:33, :487:35
      wire _T_30898 = T_23706_15 & |(io_brinfo_mask & T_26182_15_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_30900 = _T_29369 & _T_30898;	// rob.scala:484:56
      wire _T_119 = _T_30900 | _T_56 & _T_23;	// rob.scala:357:33, :487:35
      wire _T_31000 = T_23706_16 & |(io_brinfo_mask & T_26182_16_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31002 = _T_29369 & _T_31000;	// rob.scala:484:56
      wire _T_120 = _T_31002 | _T_56 & _T_24;	// rob.scala:357:33, :487:35
      wire _T_31102 = T_23706_17 & |(io_brinfo_mask & T_26182_17_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31104 = _T_29369 & _T_31102;	// rob.scala:484:56
      wire _T_121 = _T_31104 | _T_56 & _T_25;	// rob.scala:357:33, :487:35
      wire _T_31204 = T_23706_18 & |(io_brinfo_mask & T_26182_18_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31206 = _T_29369 & _T_31204;	// rob.scala:484:56
      wire _T_122 = _T_31206 | _T_56 & _T_26;	// rob.scala:357:33, :487:35
      wire _T_31306 = T_23706_19 & |(io_brinfo_mask & T_26182_19_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31308 = _T_29369 & _T_31306;	// rob.scala:484:56
      wire _T_123 = _T_31308 | _T_56 & _T_27;	// rob.scala:357:33, :487:35
      wire _T_31408 = T_23706_20 & |(io_brinfo_mask & T_26182_20_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31410 = _T_29369 & _T_31408;	// rob.scala:484:56
      wire _T_124 = _T_31410 | _T_56 & _T_28;	// rob.scala:357:33, :487:35
      wire _T_31510 = T_23706_21 & |(io_brinfo_mask & T_26182_21_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31512 = _T_29369 & _T_31510;	// rob.scala:484:56
      wire _T_125 = _T_31512 | _T_56 & _T_29;	// rob.scala:357:33, :487:35
      wire _T_31612 = T_23706_22 & |(io_brinfo_mask & T_26182_22_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31614 = _T_29369 & _T_31612;	// rob.scala:484:56
      wire _T_126 = _T_31614 | _T_56 & _T_30;	// rob.scala:357:33, :487:35
      wire _T_31714 = T_23706_23 & |(io_brinfo_mask & T_26182_23_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_31716 = _T_29369 & _T_31714;	// rob.scala:484:56
      wire _T_127 = _T_31716 | _T_56 & _T_31;	// rob.scala:357:33, :487:35
      wire _T_32082 = ~_T_3 & _T_29097;	// rob.scala:514:7, :518:7
      wire _T_32171 = io_debug_wb_valids_0 & ~_T_28590;	// rob.scala:331:55, :529:38
      wire _T_128 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, rob.scala:531:53
      wire _T_129 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h1;	// rob.scala:347:34, :531:53
      wire _T_130 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h2;	// rob.scala:347:34, :531:53
      wire _T_131 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h3;	// rob.scala:347:34, :531:53
      wire _T_132 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h4;	// rob.scala:347:34, :531:53
      wire _T_133 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h5;	// rob.scala:347:34, :531:53
      wire _T_134 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h6;	// rob.scala:347:34, :531:53
      wire _T_135 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h7;	// rob.scala:347:34, :531:53
      wire _T_136 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h8;	// rob.scala:347:34, :531:53
      wire _T_137 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h9;	// rob.scala:347:34, :531:53
      wire _T_138 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hA;	// rob.scala:347:34, :531:53
      wire _T_139 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hB;	// rob.scala:347:34, :531:53
      wire _T_140 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hC;	// rob.scala:347:34, :531:53
      wire _T_141 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hD;	// rob.scala:347:34, :531:53
      wire _T_142 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hE;	// rob.scala:347:34, :531:53
      wire _T_143 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'hF;	// rob.scala:347:34, :531:53
      wire _T_144 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h10;	// rob.scala:347:34, :531:53
      wire _T_145 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h11;	// rob.scala:347:34, :531:53
      wire _T_146 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h12;	// rob.scala:347:34, :531:53
      wire _T_147 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h13;	// rob.scala:347:34, :531:53
      wire _T_148 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h14;	// rob.scala:347:34, :531:53
      wire _T_149 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h15;	// rob.scala:347:34, :531:53
      wire _T_150 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h16;	// rob.scala:347:34, :531:53
      wire _T_151 = _io_wb_resps_0_bits_uop_rob_idx_5to1 == 5'h17;	// rob.scala:347:34, :531:53
      wire _T_32375 = io_debug_wb_valids_1 & ~_T_28598;	// rob.scala:331:55, :529:38
      wire _T_152 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, rob.scala:531:53
      wire _T_153 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h1;	// rob.scala:347:34, :531:53
      wire _T_154 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h2;	// rob.scala:347:34, :531:53
      wire _T_155 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h3;	// rob.scala:347:34, :531:53
      wire _T_156 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h4;	// rob.scala:347:34, :531:53
      wire _T_157 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h5;	// rob.scala:347:34, :531:53
      wire _T_158 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h6;	// rob.scala:347:34, :531:53
      wire _T_159 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h7;	// rob.scala:347:34, :531:53
      wire _T_160 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h8;	// rob.scala:347:34, :531:53
      wire _T_161 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h9;	// rob.scala:347:34, :531:53
      wire _T_162 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hA;	// rob.scala:347:34, :531:53
      wire _T_163 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hB;	// rob.scala:347:34, :531:53
      wire _T_164 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hC;	// rob.scala:347:34, :531:53
      wire _T_165 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hD;	// rob.scala:347:34, :531:53
      wire _T_166 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hE;	// rob.scala:347:34, :531:53
      wire _T_167 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'hF;	// rob.scala:347:34, :531:53
      wire _T_168 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h10;	// rob.scala:347:34, :531:53
      wire _T_169 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h11;	// rob.scala:347:34, :531:53
      wire _T_170 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h12;	// rob.scala:347:34, :531:53
      wire _T_171 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h13;	// rob.scala:347:34, :531:53
      wire _T_172 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h14;	// rob.scala:347:34, :531:53
      wire _T_173 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h15;	// rob.scala:347:34, :531:53
      wire _T_174 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h16;	// rob.scala:347:34, :531:53
      wire _T_175 = _io_wb_resps_1_bits_uop_rob_idx_5to1 == 5'h17;	// rob.scala:347:34, :531:53
      wire _T_32579 = io_debug_wb_valids_2 & ~_T_28606;	// rob.scala:331:55, :529:38
      wire _T_176 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, rob.scala:531:53
      wire _T_177 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h1;	// rob.scala:347:34, :531:53
      wire _T_178 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h2;	// rob.scala:347:34, :531:53
      wire _T_179 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h3;	// rob.scala:347:34, :531:53
      wire _T_180 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h4;	// rob.scala:347:34, :531:53
      wire _T_181 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h5;	// rob.scala:347:34, :531:53
      wire _T_182 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h6;	// rob.scala:347:34, :531:53
      wire _T_183 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h7;	// rob.scala:347:34, :531:53
      wire _T_184 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h8;	// rob.scala:347:34, :531:53
      wire _T_185 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h9;	// rob.scala:347:34, :531:53
      wire _T_186 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hA;	// rob.scala:347:34, :531:53
      wire _T_187 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hB;	// rob.scala:347:34, :531:53
      wire _T_188 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hC;	// rob.scala:347:34, :531:53
      wire _T_189 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hD;	// rob.scala:347:34, :531:53
      wire _T_190 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hE;	// rob.scala:347:34, :531:53
      wire _T_191 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'hF;	// rob.scala:347:34, :531:53
      wire _T_192 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h10;	// rob.scala:347:34, :531:53
      wire _T_193 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h11;	// rob.scala:347:34, :531:53
      wire _T_194 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h12;	// rob.scala:347:34, :531:53
      wire _T_195 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h13;	// rob.scala:347:34, :531:53
      wire _T_196 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h14;	// rob.scala:347:34, :531:53
      wire _T_197 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h15;	// rob.scala:347:34, :531:53
      wire _T_198 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h16;	// rob.scala:347:34, :531:53
      wire _T_199 = _io_wb_resps_2_bits_uop_rob_idx_5to1 == 5'h17;	// rob.scala:347:34, :531:53
      wire [31:0] _T_200 = ~io_dis_valids_1 | |rob_tail ? T_38110_0_inst : io_dis_uops_1_inst;	// rob.scala:192:32, :347:34, :350:34
      wire [31:0] _T_201 = io_dis_valids_1 & _T_9 ? io_dis_uops_1_inst : T_38110_1_inst;	// rob.scala:350:34
      wire [31:0] _T_202 = io_dis_valids_1 & _T_10 ? io_dis_uops_1_inst : T_38110_2_inst;	// rob.scala:350:34
      wire [31:0] _T_203 = io_dis_valids_1 & _T_11 ? io_dis_uops_1_inst : T_38110_3_inst;	// rob.scala:350:34
      wire [31:0] _T_204 = io_dis_valids_1 & _T_12 ? io_dis_uops_1_inst : T_38110_4_inst;	// rob.scala:350:34
      wire [31:0] _T_205 = io_dis_valids_1 & _T_13 ? io_dis_uops_1_inst : T_38110_5_inst;	// rob.scala:350:34
      wire [31:0] _T_206 = io_dis_valids_1 & _T_14 ? io_dis_uops_1_inst : T_38110_6_inst;	// rob.scala:350:34
      wire [31:0] _T_207 = io_dis_valids_1 & _T_15 ? io_dis_uops_1_inst : T_38110_7_inst;	// rob.scala:350:34
      wire [31:0] _T_208 = io_dis_valids_1 & _T_16 ? io_dis_uops_1_inst : T_38110_8_inst;	// rob.scala:350:34
      wire [31:0] _T_209 = io_dis_valids_1 & _T_17 ? io_dis_uops_1_inst : T_38110_9_inst;	// rob.scala:350:34
      wire [31:0] _T_210 = io_dis_valids_1 & _T_18 ? io_dis_uops_1_inst : T_38110_10_inst;	// rob.scala:350:34
      wire [31:0] _T_211 = io_dis_valids_1 & _T_19 ? io_dis_uops_1_inst : T_38110_11_inst;	// rob.scala:350:34
      wire [31:0] _T_212 = io_dis_valids_1 & _T_20 ? io_dis_uops_1_inst : T_38110_12_inst;	// rob.scala:350:34
      wire [31:0] _T_213 = io_dis_valids_1 & _T_21 ? io_dis_uops_1_inst : T_38110_13_inst;	// rob.scala:350:34
      wire [31:0] _T_214 = io_dis_valids_1 & _T_22 ? io_dis_uops_1_inst : T_38110_14_inst;	// rob.scala:350:34
      wire [31:0] _T_215 = io_dis_valids_1 & _T_23 ? io_dis_uops_1_inst : T_38110_15_inst;	// rob.scala:350:34
      wire [31:0] _T_216 = io_dis_valids_1 & _T_24 ? io_dis_uops_1_inst : T_38110_16_inst;	// rob.scala:350:34
      wire [31:0] _T_217 = io_dis_valids_1 & _T_25 ? io_dis_uops_1_inst : T_38110_17_inst;	// rob.scala:350:34
      wire [31:0] _T_218 = io_dis_valids_1 & _T_26 ? io_dis_uops_1_inst : T_38110_18_inst;	// rob.scala:350:34
      wire [31:0] _T_219 = io_dis_valids_1 & _T_27 ? io_dis_uops_1_inst : T_38110_19_inst;	// rob.scala:350:34
      wire [31:0] _T_220 = io_dis_valids_1 & _T_28 ? io_dis_uops_1_inst : T_38110_20_inst;	// rob.scala:350:34
      wire [31:0] _T_221 = io_dis_valids_1 & _T_29 ? io_dis_uops_1_inst : T_38110_21_inst;	// rob.scala:350:34
      wire [31:0] _T_222 = io_dis_valids_1 & _T_30 ? io_dis_uops_1_inst : T_38110_22_inst;	// rob.scala:350:34
      wire [31:0] _T_223 = io_dis_valids_1 & _T_31 ? io_dis_uops_1_inst : T_38110_23_inst;	// rob.scala:350:34
      wire _T_224 = ~io_dis_valids_1 & _T_23559 & ~casez_tmp_93;	// rob.scala:346:7, :355:47, :356:7
      wire _T_40551 = io_brinfo_valid & _T_28620;	// rob.scala:400:29
      wire _T_41296 = T_35634_0 & |(io_brinfo_mask & T_38110_0_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41298 = _T_29369 & _T_41296;	// rob.scala:484:56
      wire _T_225 = _T_41298 | ~(~_T_224 | |rob_tail);	// rob.scala:192:32, :347:34, :357:33, :487:35
      wire _T_41398 = T_35634_1 & |(io_brinfo_mask & T_38110_1_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41400 = _T_29369 & _T_41398;	// rob.scala:484:56
      wire _T_226 = _T_41400 | _T_224 & _T_9;	// rob.scala:357:33, :487:35
      wire _T_41500 = T_35634_2 & |(io_brinfo_mask & T_38110_2_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41502 = _T_29369 & _T_41500;	// rob.scala:484:56
      wire _T_227 = _T_41502 | _T_224 & _T_10;	// rob.scala:357:33, :487:35
      wire _T_41602 = T_35634_3 & |(io_brinfo_mask & T_38110_3_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41604 = _T_29369 & _T_41602;	// rob.scala:484:56
      wire _T_228 = _T_41604 | _T_224 & _T_11;	// rob.scala:357:33, :487:35
      wire _T_41704 = T_35634_4 & |(io_brinfo_mask & T_38110_4_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41706 = _T_29369 & _T_41704;	// rob.scala:484:56
      wire _T_229 = _T_41706 | _T_224 & _T_12;	// rob.scala:357:33, :487:35
      wire _T_41806 = T_35634_5 & |(io_brinfo_mask & T_38110_5_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41808 = _T_29369 & _T_41806;	// rob.scala:484:56
      wire _T_230 = _T_41808 | _T_224 & _T_13;	// rob.scala:357:33, :487:35
      wire _T_41908 = T_35634_6 & |(io_brinfo_mask & T_38110_6_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_41910 = _T_29369 & _T_41908;	// rob.scala:484:56
      wire _T_231 = _T_41910 | _T_224 & _T_14;	// rob.scala:357:33, :487:35
      wire _T_42010 = T_35634_7 & |(io_brinfo_mask & T_38110_7_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42012 = _T_29369 & _T_42010;	// rob.scala:484:56
      wire _T_232 = _T_42012 | _T_224 & _T_15;	// rob.scala:357:33, :487:35
      wire _T_42112 = T_35634_8 & |(io_brinfo_mask & T_38110_8_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42114 = _T_29369 & _T_42112;	// rob.scala:484:56
      wire _T_233 = _T_42114 | _T_224 & _T_16;	// rob.scala:357:33, :487:35
      wire _T_42214 = T_35634_9 & |(io_brinfo_mask & T_38110_9_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42216 = _T_29369 & _T_42214;	// rob.scala:484:56
      wire _T_234 = _T_42216 | _T_224 & _T_17;	// rob.scala:357:33, :487:35
      wire _T_42316 = T_35634_10 & |(io_brinfo_mask & T_38110_10_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42318 = _T_29369 & _T_42316;	// rob.scala:484:56
      wire _T_235 = _T_42318 | _T_224 & _T_18;	// rob.scala:357:33, :487:35
      wire _T_42418 = T_35634_11 & |(io_brinfo_mask & T_38110_11_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42420 = _T_29369 & _T_42418;	// rob.scala:484:56
      wire _T_236 = _T_42420 | _T_224 & _T_19;	// rob.scala:357:33, :487:35
      wire _T_42520 = T_35634_12 & |(io_brinfo_mask & T_38110_12_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42522 = _T_29369 & _T_42520;	// rob.scala:484:56
      wire _T_237 = _T_42522 | _T_224 & _T_20;	// rob.scala:357:33, :487:35
      wire _T_42622 = T_35634_13 & |(io_brinfo_mask & T_38110_13_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42624 = _T_29369 & _T_42622;	// rob.scala:484:56
      wire _T_238 = _T_42624 | _T_224 & _T_21;	// rob.scala:357:33, :487:35
      wire _T_42724 = T_35634_14 & |(io_brinfo_mask & T_38110_14_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42726 = _T_29369 & _T_42724;	// rob.scala:484:56
      wire _T_239 = _T_42726 | _T_224 & _T_22;	// rob.scala:357:33, :487:35
      wire _T_42826 = T_35634_15 & |(io_brinfo_mask & T_38110_15_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42828 = _T_29369 & _T_42826;	// rob.scala:484:56
      wire _T_240 = _T_42828 | _T_224 & _T_23;	// rob.scala:357:33, :487:35
      wire _T_42928 = T_35634_16 & |(io_brinfo_mask & T_38110_16_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_42930 = _T_29369 & _T_42928;	// rob.scala:484:56
      wire _T_241 = _T_42930 | _T_224 & _T_24;	// rob.scala:357:33, :487:35
      wire _T_43030 = T_35634_17 & |(io_brinfo_mask & T_38110_17_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43032 = _T_29369 & _T_43030;	// rob.scala:484:56
      wire _T_242 = _T_43032 | _T_224 & _T_25;	// rob.scala:357:33, :487:35
      wire _T_43132 = T_35634_18 & |(io_brinfo_mask & T_38110_18_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43134 = _T_29369 & _T_43132;	// rob.scala:484:56
      wire _T_243 = _T_43134 | _T_224 & _T_26;	// rob.scala:357:33, :487:35
      wire _T_43234 = T_35634_19 & |(io_brinfo_mask & T_38110_19_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43236 = _T_29369 & _T_43234;	// rob.scala:484:56
      wire _T_244 = _T_43236 | _T_224 & _T_27;	// rob.scala:357:33, :487:35
      wire _T_43336 = T_35634_20 & |(io_brinfo_mask & T_38110_20_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43338 = _T_29369 & _T_43336;	// rob.scala:484:56
      wire _T_245 = _T_43338 | _T_224 & _T_28;	// rob.scala:357:33, :487:35
      wire _T_43438 = T_35634_21 & |(io_brinfo_mask & T_38110_21_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43440 = _T_29369 & _T_43438;	// rob.scala:484:56
      wire _T_246 = _T_43440 | _T_224 & _T_29;	// rob.scala:357:33, :487:35
      wire _T_43540 = T_35634_22 & |(io_brinfo_mask & T_38110_22_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43542 = _T_29369 & _T_43540;	// rob.scala:484:56
      wire _T_247 = _T_43542 | _T_224 & _T_30;	// rob.scala:357:33, :487:35
      wire _T_43642 = T_35634_23 & |(io_brinfo_mask & T_38110_23_br_mask);	// rob.scala:347:34, :350:34, :481:39, util.scala:45:{52,60}
      wire _T_43644 = _T_29369 & _T_43642;	// rob.scala:484:56
      wire _T_248 = _T_43644 | _T_224 & _T_31;	// rob.scala:357:33, :487:35
      wire _T_44010 = ~_T_4 & _T_29097;	// rob.scala:514:7, :518:7
      wire _T_44099 = io_debug_wb_valids_0 & _T_28590;	// rob.scala:529:38
      wire _T_44303 = io_debug_wb_valids_1 & _T_28598;	// rob.scala:529:38
      wire _T_44507 = io_debug_wb_valids_2 & _T_28606;	// rob.scala:529:38
      wire _T_47869 = io_dis_valids_0 & io_dis_uops_0_exception;	// rob.scala:656:40
      wire _T_47875 = ~(T_47616 | _T_47568) & rob_state != 2'h2;	// rob.scala:443:23, :612:22, :659:{10,30,51,64}
      wire _T_47876 = io_lxcpt_valid | io_bxcpt_valid;	// rob.scala:661:28
      wire _T_47887 = io_lxcpt_valid & ~io_bxcpt_valid | io_lxcpt_valid & io_bxcpt_valid &
                {io_lxcpt_bits_uop_rob_idx <= _rob_tail_idx, io_lxcpt_bits_uop_rob_idx} <
                {io_bxcpt_bits_uop_rob_idx <= _rob_tail_idx, io_bxcpt_bits_uop_rob_idx};	// Cat.scala:20:58, rob.scala:650:{58,71,80}, :663:{46,49,66}, :664:64
      wire [5:0] _T_47888_rob_idx = _T_47887 ? io_lxcpt_bits_uop_rob_idx : io_bxcpt_bits_uop_rob_idx;	// rob.scala:666:32
      wire _T_47981 = ~r_xcpt_val | {_T_47888_rob_idx <= _rob_tail_idx, _T_47888_rob_idx} < {r_xcpt_uop_rob_idx
                <= _rob_tail_idx, r_xcpt_uop_rob_idx};	// Cat.scala:20:58, rob.scala:650:{58,71,80}, :667:{16,28}
      wire _T_249 = ~_T_47876 & ~r_xcpt_val & (_T_47869 | io_dis_valids_1 & io_dis_uops_1_exception);	// rob.scala:656:40, :662:7, :667:16, :675:{18,51}, :676:7
      wire [7:0] _T_250 = _T_47875 ? (_T_249 ? (_T_47869 ? io_dis_uops_0_br_mask : io_dis_uops_1_br_mask) : _T_47876
                & _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_br_mask : io_bxcpt_bits_uop_br_mask) :
                r_xcpt_uop_br_mask) : r_xcpt_uop_br_mask;	// rob.scala:666:32, :670:37, :681:26
  always @(posedge clk) begin	// rob.scala:350:34
    if (reset) begin	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      rob_state <= 2'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:{5,59}
      rob_head <= 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:{5,58}
      rob_tail <= 5'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, :14:5
      r_xcpt_val <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :36:5
      r_partial_row <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :125:5
      T_23706_0 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_1 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_2 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_3 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_4 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_5 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_6 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_7 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_8 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_9 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_10 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_11 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_12 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_13 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_14 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_15 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_16 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_17 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_18 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_19 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_20 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_21 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_22 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_23706_23 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :187:5
      T_35634_0 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_1 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_2 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_3 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_4 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_5 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_6 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_7 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_8 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_9 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_10 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_11 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_12 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_13 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_14 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_15 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_16 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_17 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_18 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_19 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_20 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_21 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_22 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
      T_35634_23 <= 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :1555:5
    end
    else begin	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:5
      r_partial_row <= ~_T_23652 & _T_23559 & ~io_dis_new_packet | _T_23652 ? io_dis_partial_stall : r_partial_row;	// rob.scala:298:4, :301:21, :303:44, :304:4, :305:21
      T_23706_0 <= (~_T_3 | |rob_head) & ~_T_29370 & (~_T_29097 | |_T_2) & (io_dis_valids_0 & ~(|rob_tail) |
                                                T_23706_0);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :347:34, :459:33, :486:24, :500:28
      T_23706_1 <= (~_T_3 | ~_T_81) & ~_T_29472 & (~_T_29097 | _T_2 != 5'h1) & (io_dis_valids_0 & _T_9 |
                                                T_23706_1);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_2 <= (~_T_3 | ~_T_82) & ~_T_29574 & (~_T_29097 | _T_2 != 5'h2) & (io_dis_valids_0 & _T_10 |
                                                T_23706_2);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_3 <= (~_T_3 | ~_T_83) & ~_T_29676 & (~_T_29097 | _T_2 != 5'h3) & (io_dis_valids_0 & _T_11 |
                                                T_23706_3);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_4 <= (~_T_3 | ~_T_84) & ~_T_29778 & (~_T_29097 | _T_2 != 5'h4) & (io_dis_valids_0 & _T_12 |
                                                T_23706_4);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_5 <= (~_T_3 | ~_T_85) & ~_T_29880 & (~_T_29097 | _T_2 != 5'h5) & (io_dis_valids_0 & _T_13 |
                                                T_23706_5);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_6 <= (~_T_3 | ~_T_86) & ~_T_29982 & (~_T_29097 | _T_2 != 5'h6) & (io_dis_valids_0 & _T_14 |
                                                T_23706_6);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_7 <= (~_T_3 | ~_T_87) & ~_T_30084 & (~_T_29097 | _T_2 != 5'h7) & (io_dis_valids_0 & _T_15 |
                                                T_23706_7);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_8 <= (~_T_3 | ~_T_88) & ~_T_30186 & (~_T_29097 | _T_2 != 5'h8) & (io_dis_valids_0 & _T_16 |
                                                T_23706_8);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_9 <= (~_T_3 | ~_T_89) & ~_T_30288 & (~_T_29097 | _T_2 != 5'h9) & (io_dis_valids_0 & _T_17 |
                                                T_23706_9);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_10 <= (~_T_3 | ~_T_90) & ~_T_30390 & (~_T_29097 | _T_2 != 5'hA) & (io_dis_valids_0 & _T_18 |
                                                T_23706_10);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_11 <= (~_T_3 | ~_T_91) & ~_T_30492 & (~_T_29097 | _T_2 != 5'hB) & (io_dis_valids_0 & _T_19 |
                                                T_23706_11);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_12 <= (~_T_3 | ~_T_92) & ~_T_30594 & (~_T_29097 | _T_2 != 5'hC) & (io_dis_valids_0 & _T_20 |
                                                T_23706_12);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_13 <= (~_T_3 | ~_T_93) & ~_T_30696 & (~_T_29097 | _T_2 != 5'hD) & (io_dis_valids_0 & _T_21 |
                                                T_23706_13);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_14 <= (~_T_3 | ~_T_94) & ~_T_30798 & (~_T_29097 | _T_2 != 5'hE) & (io_dis_valids_0 & _T_22 |
                                                T_23706_14);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_15 <= (~_T_3 | ~_T_95) & ~_T_30900 & (~_T_29097 | _T_2 != 5'hF) & (io_dis_valids_0 & _T_23 |
                                                T_23706_15);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_16 <= (~_T_3 | ~_T_96) & ~_T_31002 & (~_T_29097 | _T_2 != 5'h10) & (io_dis_valids_0 & _T_24 |
                                                T_23706_16);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_17 <= (~_T_3 | ~_T_97) & ~_T_31104 & (~_T_29097 | _T_2 != 5'h11) & (io_dis_valids_0 & _T_25 |
                                                T_23706_17);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_18 <= (~_T_3 | ~_T_98) & ~_T_31206 & (~_T_29097 | _T_2 != 5'h12) & (io_dis_valids_0 & _T_26 |
                                                T_23706_18);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_19 <= (~_T_3 | ~_T_99) & ~_T_31308 & (~_T_29097 | _T_2 != 5'h13) & (io_dis_valids_0 & _T_27 |
                                                T_23706_19);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_20 <= (~_T_3 | ~_T_100) & ~_T_31410 & (~_T_29097 | _T_2 != 5'h14) & (io_dis_valids_0 & _T_28 |
                                                T_23706_20);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_21 <= (~_T_3 | ~_T_101) & ~_T_31512 & (~_T_29097 | _T_2 != 5'h15) & (io_dis_valids_0 & _T_29 |
                                                T_23706_21);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_22 <= (~_T_3 | ~_T_102) & ~_T_31614 & (~_T_29097 | _T_2 != 5'h16) & (io_dis_valids_0 & _T_30 |
                                                T_23706_22);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_23706_23 <= (~_T_3 | ~_T_103) & ~_T_31716 & (~_T_29097 | _T_2 != 5'h17) & (io_dis_valids_0 & _T_31 |
                                                T_23706_23);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_0 <= (~_T_4 | |rob_head) & ~_T_41298 & (~_T_29097 | |_T_2) & (io_dis_valids_1 & ~(|rob_tail) |
                                                T_35634_0);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :347:34, :459:33, :486:24, :500:28
      T_35634_1 <= (~_T_4 | ~_T_81) & ~_T_41400 & (~_T_29097 | _T_2 != 5'h1) & (io_dis_valids_1 & _T_9 |
                                                T_35634_1);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_2 <= (~_T_4 | ~_T_82) & ~_T_41502 & (~_T_29097 | _T_2 != 5'h2) & (io_dis_valids_1 & _T_10 |
                                                T_35634_2);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_3 <= (~_T_4 | ~_T_83) & ~_T_41604 & (~_T_29097 | _T_2 != 5'h3) & (io_dis_valids_1 & _T_11 |
                                                T_35634_3);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_4 <= (~_T_4 | ~_T_84) & ~_T_41706 & (~_T_29097 | _T_2 != 5'h4) & (io_dis_valids_1 & _T_12 |
                                                T_35634_4);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_5 <= (~_T_4 | ~_T_85) & ~_T_41808 & (~_T_29097 | _T_2 != 5'h5) & (io_dis_valids_1 & _T_13 |
                                                T_35634_5);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_6 <= (~_T_4 | ~_T_86) & ~_T_41910 & (~_T_29097 | _T_2 != 5'h6) & (io_dis_valids_1 & _T_14 |
                                                T_35634_6);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_7 <= (~_T_4 | ~_T_87) & ~_T_42012 & (~_T_29097 | _T_2 != 5'h7) & (io_dis_valids_1 & _T_15 |
                                                T_35634_7);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_8 <= (~_T_4 | ~_T_88) & ~_T_42114 & (~_T_29097 | _T_2 != 5'h8) & (io_dis_valids_1 & _T_16 |
                                                T_35634_8);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_9 <= (~_T_4 | ~_T_89) & ~_T_42216 & (~_T_29097 | _T_2 != 5'h9) & (io_dis_valids_1 & _T_17 |
                                                T_35634_9);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_10 <= (~_T_4 | ~_T_90) & ~_T_42318 & (~_T_29097 | _T_2 != 5'hA) & (io_dis_valids_1 & _T_18 |
                                                T_35634_10);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_11 <= (~_T_4 | ~_T_91) & ~_T_42420 & (~_T_29097 | _T_2 != 5'hB) & (io_dis_valids_1 & _T_19 |
                                                T_35634_11);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_12 <= (~_T_4 | ~_T_92) & ~_T_42522 & (~_T_29097 | _T_2 != 5'hC) & (io_dis_valids_1 & _T_20 |
                                                T_35634_12);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_13 <= (~_T_4 | ~_T_93) & ~_T_42624 & (~_T_29097 | _T_2 != 5'hD) & (io_dis_valids_1 & _T_21 |
                                                T_35634_13);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_14 <= (~_T_4 | ~_T_94) & ~_T_42726 & (~_T_29097 | _T_2 != 5'hE) & (io_dis_valids_1 & _T_22 |
                                                T_35634_14);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_15 <= (~_T_4 | ~_T_95) & ~_T_42828 & (~_T_29097 | _T_2 != 5'hF) & (io_dis_valids_1 & _T_23 |
                                                T_35634_15);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_16 <= (~_T_4 | ~_T_96) & ~_T_42930 & (~_T_29097 | _T_2 != 5'h10) & (io_dis_valids_1 & _T_24 |
                                                T_35634_16);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_17 <= (~_T_4 | ~_T_97) & ~_T_43032 & (~_T_29097 | _T_2 != 5'h11) & (io_dis_valids_1 & _T_25 |
                                                T_35634_17);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_18 <= (~_T_4 | ~_T_98) & ~_T_43134 & (~_T_29097 | _T_2 != 5'h12) & (io_dis_valids_1 & _T_26 |
                                                T_35634_18);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_19 <= (~_T_4 | ~_T_99) & ~_T_43236 & (~_T_29097 | _T_2 != 5'h13) & (io_dis_valids_1 & _T_27 |
                                                T_35634_19);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_20 <= (~_T_4 | ~_T_100) & ~_T_43338 & (~_T_29097 | _T_2 != 5'h14) & (io_dis_valids_1 & _T_28 |
                                                T_35634_20);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_21 <= (~_T_4 | ~_T_101) & ~_T_43440 & (~_T_29097 | _T_2 != 5'h15) & (io_dis_valids_1 & _T_29 |
                                                T_35634_21);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_22 <= (~_T_4 | ~_T_102) & ~_T_43542 & (~_T_29097 | _T_2 != 5'h16) & (io_dis_valids_1 & _T_30 |
                                                T_35634_22);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      T_35634_23 <= (~_T_4 | ~_T_103) & ~_T_43644 & (~_T_29097 | _T_2 != 5'h17) & (io_dis_valids_1 & _T_31 |
                                                T_35634_23);	// rob.scala:347:34, :451:58, :459:33, :486:24, :500:28
      r_xcpt_val <= ~(T_47616 | _T_29369 & |(io_brinfo_mask & _T_250)) & (_T_47875 & (_T_249 | _T_47876 &
                                                _T_47981) | r_xcpt_val);	// rob.scala:612:22, :667:16, :669:37, :680:26, :688:28, :690:18, util.scala:23:33, :45:{52,60}
      rob_head <= _T ? (rob_head == 5'h17 ? 5'h0 : rob_head + 5'h1) : rob_head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, :149:5, rob.scala:347:34, :716:89, :720:16, util.scala:75:28, :76:{13,35}
      rob_tail <= ~_T_48144 & ~_T_29369 & |{io_dis_valids_1, io_dis_valids_0} & ~io_dis_partial_stall ?
                                                (rob_tail == 5'h17 ? 5'h0 : rob_tail + 5'h1) : ~_T_48144 & _T_29369 ?
                                                (_io_brinfo_rob_idx_5to1 == 5'h17 ? 5'h0 : _io_brinfo_rob_idx_5to1 + 5'h1) : _T_48144 ?
                                                (|rob_tail ? rob_tail - 5'h1 : 5'h17) : rob_tail;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58, :104:20, rob.scala:192:32, :347:34, :727:4, :728:16, :731:4, :732:16, :734:{36,51}, :735:4, :736:16, util.scala:75:28, :76:{13,35}, :92:{13,39}
      rob_state <= &rob_state ? (~_T_47568 & _T_48195 ? 2'h1 : _T_47568 ? 2'h2 : _T_8) : _T_8;	// Conditional.scala:24:42, rob.scala:443:23, :453:100, :806:13, :807:26, :810:13, :811:26
    end
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (~(~io_dis_valids_0 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_26182_0_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_9)	// rob.scala:350:34
      T_26182_1_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_10)	// rob.scala:350:34
      T_26182_2_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_11)	// rob.scala:350:34
      T_26182_3_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_12)	// rob.scala:350:34
      T_26182_4_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_13)	// rob.scala:350:34
      T_26182_5_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_14)	// rob.scala:350:34
      T_26182_6_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_15)	// rob.scala:350:34
      T_26182_7_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_16)	// rob.scala:350:34
      T_26182_8_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_17)	// rob.scala:350:34
      T_26182_9_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_18)	// rob.scala:350:34
      T_26182_10_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_19)	// rob.scala:350:34
      T_26182_11_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_20)	// rob.scala:350:34
      T_26182_12_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_21)	// rob.scala:350:34
      T_26182_13_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_22)	// rob.scala:350:34
      T_26182_14_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_23)	// rob.scala:350:34
      T_26182_15_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_24)	// rob.scala:350:34
      T_26182_16_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_25)	// rob.scala:350:34
      T_26182_17_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_26)	// rob.scala:350:34
      T_26182_18_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_27)	// rob.scala:350:34
      T_26182_19_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_28)	// rob.scala:350:34
      T_26182_20_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_29)	// rob.scala:350:34
      T_26182_21_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_30)	// rob.scala:350:34
      T_26182_22_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_valid <= io_dis_uops_0_valid;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_iw_state <= io_dis_uops_0_iw_state;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_uopc <= io_dis_uops_0_uopc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_pc <= io_dis_uops_0_pc;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_fu_code <= io_dis_uops_0_fu_code;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_br_type <= io_dis_uops_0_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_op1_sel <= io_dis_uops_0_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_op2_sel <= io_dis_uops_0_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_imm_sel <= io_dis_uops_0_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_op_fcn <= io_dis_uops_0_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_fcn_dw <= io_dis_uops_0_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_rf_wen <= io_dis_uops_0_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_csr_cmd <= io_dis_uops_0_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_is_load <= io_dis_uops_0_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_is_sta <= io_dis_uops_0_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ctrl_is_std <= io_dis_uops_0_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_wakeup_delay <= io_dis_uops_0_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_allocate_brtag <= io_dis_uops_0_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_br_or_jmp <= io_dis_uops_0_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_jump <= io_dis_uops_0_is_jump;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_jal <= io_dis_uops_0_is_jal;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_ret <= io_dis_uops_0_is_ret;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_call <= io_dis_uops_0_is_call;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_tag <= io_dis_uops_0_br_tag;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_prediction_bpd_predict_val <= io_dis_uops_0_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_prediction_bpd_predict_taken <= io_dis_uops_0_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_prediction_btb_hit <= io_dis_uops_0_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_prediction_btb_predicted <= io_dis_uops_0_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_br_prediction_is_br_or_jalr <= io_dis_uops_0_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_fetch_pc_lob <= io_dis_uops_0_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_imm_packed <= io_dis_uops_0_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_csr_addr <= io_dis_uops_0_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_rob_idx <= io_dis_uops_0_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ldq_idx <= io_dis_uops_0_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_stq_idx <= io_dis_uops_0_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_brob_idx <= io_dis_uops_0_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_pdst <= io_dis_uops_0_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_pop1 <= io_dis_uops_0_pop1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_pop2 <= io_dis_uops_0_pop2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_pop3 <= io_dis_uops_0_pop3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_prs1_busy <= io_dis_uops_0_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_prs2_busy <= io_dis_uops_0_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_prs3_busy <= io_dis_uops_0_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_stale_pdst <= io_dis_uops_0_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_exception <= io_dis_uops_0_exception;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_exc_cause <= io_dis_uops_0_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_bypassable <= io_dis_uops_0_bypassable;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_mem_cmd <= io_dis_uops_0_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_mem_typ <= io_dis_uops_0_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_fence <= io_dis_uops_0_is_fence;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_fencei <= io_dis_uops_0_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_store <= io_dis_uops_0_is_store;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_amo <= io_dis_uops_0_is_amo;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_load <= io_dis_uops_0_is_load;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_is_unique <= io_dis_uops_0_is_unique;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_flush_on_commit <= io_dis_uops_0_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ldst <= io_dis_uops_0_ldst;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_lrs1 <= io_dis_uops_0_lrs1;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_lrs2 <= io_dis_uops_0_lrs2;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_lrs3 <= io_dis_uops_0_lrs3;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_ldst_val <= io_dis_uops_0_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_dst_rtype <= io_dis_uops_0_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_lrs1_rtype <= io_dis_uops_0_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_lrs2_rtype <= io_dis_uops_0_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_frs3_en <= io_dis_uops_0_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_fp_val <= io_dis_uops_0_fp_val;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_fp_single <= io_dis_uops_0_fp_single;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_xcpt_if <= io_dis_uops_0_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_replay_if <= io_dis_uops_0_replay_if;	// rob.scala:350:34
    if (io_dis_valids_0 & _T_31)	// rob.scala:350:34
      T_26182_23_debug_events_fetch_seq <= io_dis_uops_0_debug_events_fetch_seq;	// rob.scala:350:34
    T_26182_0_stat_brjmp_mispredicted <= _T_28623 & _T_57 ? io_brinfo_mispredict : io_dis_valids_0 ? |rob_tail & (|rob_tail ?
                                T_26182_0_stat_brjmp_mispredicted : io_dis_uops_0_stat_brjmp_mispredicted) :
                                T_26182_0_stat_brjmp_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :353:52, :402:72
    T_26182_1_stat_brjmp_mispredicted <= _T_28623 & _T_58 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_9 & (_T_9 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_1_stat_brjmp_mispredicted) :
                                T_26182_1_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_2_stat_brjmp_mispredicted <= _T_28623 & _T_59 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_10 & (_T_10 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_2_stat_brjmp_mispredicted) :
                                T_26182_2_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_3_stat_brjmp_mispredicted <= _T_28623 & _T_60 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_11 & (_T_11 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_3_stat_brjmp_mispredicted) :
                                T_26182_3_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_4_stat_brjmp_mispredicted <= _T_28623 & _T_61 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_12 & (_T_12 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_4_stat_brjmp_mispredicted) :
                                T_26182_4_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_5_stat_brjmp_mispredicted <= _T_28623 & _T_62 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_13 & (_T_13 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_5_stat_brjmp_mispredicted) :
                                T_26182_5_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_6_stat_brjmp_mispredicted <= _T_28623 & _T_63 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_14 & (_T_14 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_6_stat_brjmp_mispredicted) :
                                T_26182_6_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_7_stat_brjmp_mispredicted <= _T_28623 & _T_64 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_15 & (_T_15 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_7_stat_brjmp_mispredicted) :
                                T_26182_7_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_8_stat_brjmp_mispredicted <= _T_28623 & _T_65 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_16 & (_T_16 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_8_stat_brjmp_mispredicted) :
                                T_26182_8_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_9_stat_brjmp_mispredicted <= _T_28623 & _T_66 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_17 & (_T_17 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_9_stat_brjmp_mispredicted) :
                                T_26182_9_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_10_stat_brjmp_mispredicted <= _T_28623 & _T_67 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_18 & (_T_18 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_10_stat_brjmp_mispredicted) :
                                T_26182_10_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_11_stat_brjmp_mispredicted <= _T_28623 & _T_68 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_19 & (_T_19 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_11_stat_brjmp_mispredicted) :
                                T_26182_11_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_12_stat_brjmp_mispredicted <= _T_28623 & _T_69 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_20 & (_T_20 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_12_stat_brjmp_mispredicted) :
                                T_26182_12_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_13_stat_brjmp_mispredicted <= _T_28623 & _T_70 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_21 & (_T_21 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_13_stat_brjmp_mispredicted) :
                                T_26182_13_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_14_stat_brjmp_mispredicted <= _T_28623 & _T_71 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_22 & (_T_22 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_14_stat_brjmp_mispredicted) :
                                T_26182_14_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_15_stat_brjmp_mispredicted <= _T_28623 & _T_72 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_23 & (_T_23 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_15_stat_brjmp_mispredicted) :
                                T_26182_15_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_16_stat_brjmp_mispredicted <= _T_28623 & _T_73 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_24 & (_T_24 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_16_stat_brjmp_mispredicted) :
                                T_26182_16_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_17_stat_brjmp_mispredicted <= _T_28623 & _T_74 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_25 & (_T_25 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_17_stat_brjmp_mispredicted) :
                                T_26182_17_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_18_stat_brjmp_mispredicted <= _T_28623 & _T_75 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_26 & (_T_26 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_18_stat_brjmp_mispredicted) :
                                T_26182_18_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_19_stat_brjmp_mispredicted <= _T_28623 & _T_76 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_27 & (_T_27 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_19_stat_brjmp_mispredicted) :
                                T_26182_19_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_20_stat_brjmp_mispredicted <= _T_28623 & _T_77 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_28 & (_T_28 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_20_stat_brjmp_mispredicted) :
                                T_26182_20_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_21_stat_brjmp_mispredicted <= _T_28623 & _T_78 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_29 & (_T_29 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_21_stat_brjmp_mispredicted) :
                                T_26182_21_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_22_stat_brjmp_mispredicted <= _T_28623 & _T_79 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_30 & (_T_30 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_22_stat_brjmp_mispredicted) :
                                T_26182_22_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_23_stat_brjmp_mispredicted <= _T_28623 & _T_80 ? io_brinfo_mispredict : io_dis_valids_0 ? ~_T_31 & (_T_31 ?
                                io_dis_uops_0_stat_brjmp_mispredicted : T_26182_23_stat_brjmp_mispredicted) :
                                T_26182_23_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_26182_0_stat_btb_mispredicted <= _T_28623 & _T_57 ? io_brinfo_btb_mispredict : ~io_dis_valids_0 | |rob_tail ?
                                T_26182_0_stat_btb_mispredicted : io_dis_uops_0_stat_btb_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :403:72
    T_26182_1_stat_btb_mispredicted <= _T_28623 & _T_58 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_9 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_1_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_2_stat_btb_mispredicted <= _T_28623 & _T_59 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_10 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_2_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_3_stat_btb_mispredicted <= _T_28623 & _T_60 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_11 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_3_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_4_stat_btb_mispredicted <= _T_28623 & _T_61 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_12 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_4_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_5_stat_btb_mispredicted <= _T_28623 & _T_62 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_13 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_5_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_6_stat_btb_mispredicted <= _T_28623 & _T_63 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_14 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_6_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_7_stat_btb_mispredicted <= _T_28623 & _T_64 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_15 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_7_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_8_stat_btb_mispredicted <= _T_28623 & _T_65 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_16 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_8_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_9_stat_btb_mispredicted <= _T_28623 & _T_66 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_17 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_9_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_10_stat_btb_mispredicted <= _T_28623 & _T_67 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_18 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_10_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_11_stat_btb_mispredicted <= _T_28623 & _T_68 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_19 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_11_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_12_stat_btb_mispredicted <= _T_28623 & _T_69 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_20 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_12_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_13_stat_btb_mispredicted <= _T_28623 & _T_70 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_21 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_13_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_14_stat_btb_mispredicted <= _T_28623 & _T_71 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_22 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_14_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_15_stat_btb_mispredicted <= _T_28623 & _T_72 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_23 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_15_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_16_stat_btb_mispredicted <= _T_28623 & _T_73 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_24 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_16_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_17_stat_btb_mispredicted <= _T_28623 & _T_74 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_25 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_17_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_18_stat_btb_mispredicted <= _T_28623 & _T_75 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_26 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_18_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_19_stat_btb_mispredicted <= _T_28623 & _T_76 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_27 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_19_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_20_stat_btb_mispredicted <= _T_28623 & _T_77 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_28 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_20_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_21_stat_btb_mispredicted <= _T_28623 & _T_78 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_29 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_21_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_22_stat_btb_mispredicted <= _T_28623 & _T_79 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_30 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_22_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_23_stat_btb_mispredicted <= _T_28623 & _T_80 ? io_brinfo_btb_mispredict : io_dis_valids_0 & _T_31 ?
                                io_dis_uops_0_stat_btb_mispredicted : T_26182_23_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_26182_0_stat_btb_made_pred <= _T_28623 & _T_57 ? io_brinfo_btb_made_pred : ~io_dis_valids_0 | |rob_tail ?
                                T_26182_0_stat_btb_made_pred : io_dis_uops_0_stat_btb_made_pred;	// rob.scala:192:32, :347:34, :350:34, :404:72
    T_26182_1_stat_btb_made_pred <= _T_28623 & _T_58 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_9 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_1_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_2_stat_btb_made_pred <= _T_28623 & _T_59 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_10 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_2_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_3_stat_btb_made_pred <= _T_28623 & _T_60 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_11 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_3_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_4_stat_btb_made_pred <= _T_28623 & _T_61 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_12 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_4_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_5_stat_btb_made_pred <= _T_28623 & _T_62 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_13 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_5_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_6_stat_btb_made_pred <= _T_28623 & _T_63 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_14 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_6_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_7_stat_btb_made_pred <= _T_28623 & _T_64 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_15 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_7_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_8_stat_btb_made_pred <= _T_28623 & _T_65 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_16 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_8_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_9_stat_btb_made_pred <= _T_28623 & _T_66 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_17 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_9_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_10_stat_btb_made_pred <= _T_28623 & _T_67 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_18 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_10_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_11_stat_btb_made_pred <= _T_28623 & _T_68 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_19 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_11_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_12_stat_btb_made_pred <= _T_28623 & _T_69 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_20 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_12_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_13_stat_btb_made_pred <= _T_28623 & _T_70 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_21 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_13_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_14_stat_btb_made_pred <= _T_28623 & _T_71 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_22 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_14_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_15_stat_btb_made_pred <= _T_28623 & _T_72 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_23 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_15_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_16_stat_btb_made_pred <= _T_28623 & _T_73 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_24 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_16_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_17_stat_btb_made_pred <= _T_28623 & _T_74 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_25 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_17_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_18_stat_btb_made_pred <= _T_28623 & _T_75 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_26 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_18_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_19_stat_btb_made_pred <= _T_28623 & _T_76 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_27 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_19_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_20_stat_btb_made_pred <= _T_28623 & _T_77 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_28 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_20_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_21_stat_btb_made_pred <= _T_28623 & _T_78 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_29 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_21_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_22_stat_btb_made_pred <= _T_28623 & _T_79 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_30 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_22_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_23_stat_btb_made_pred <= _T_28623 & _T_80 ? io_brinfo_btb_made_pred : io_dis_valids_0 & _T_31 ?
                                io_dis_uops_0_stat_btb_made_pred : T_26182_23_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_26182_0_stat_bpd_mispredicted <= _T_28623 & _T_57 ? io_brinfo_bpd_mispredict : ~io_dis_valids_0 | |rob_tail ?
                                T_26182_0_stat_bpd_mispredicted : io_dis_uops_0_stat_bpd_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :405:72
    T_26182_1_stat_bpd_mispredicted <= _T_28623 & _T_58 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_9 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_1_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_2_stat_bpd_mispredicted <= _T_28623 & _T_59 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_10 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_2_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_3_stat_bpd_mispredicted <= _T_28623 & _T_60 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_11 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_3_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_4_stat_bpd_mispredicted <= _T_28623 & _T_61 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_12 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_4_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_5_stat_bpd_mispredicted <= _T_28623 & _T_62 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_13 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_5_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_6_stat_bpd_mispredicted <= _T_28623 & _T_63 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_14 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_6_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_7_stat_bpd_mispredicted <= _T_28623 & _T_64 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_15 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_7_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_8_stat_bpd_mispredicted <= _T_28623 & _T_65 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_16 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_8_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_9_stat_bpd_mispredicted <= _T_28623 & _T_66 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_17 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_9_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_10_stat_bpd_mispredicted <= _T_28623 & _T_67 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_18 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_10_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_11_stat_bpd_mispredicted <= _T_28623 & _T_68 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_19 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_11_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_12_stat_bpd_mispredicted <= _T_28623 & _T_69 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_20 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_12_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_13_stat_bpd_mispredicted <= _T_28623 & _T_70 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_21 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_13_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_14_stat_bpd_mispredicted <= _T_28623 & _T_71 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_22 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_14_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_15_stat_bpd_mispredicted <= _T_28623 & _T_72 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_23 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_15_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_16_stat_bpd_mispredicted <= _T_28623 & _T_73 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_24 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_16_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_17_stat_bpd_mispredicted <= _T_28623 & _T_74 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_25 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_17_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_18_stat_bpd_mispredicted <= _T_28623 & _T_75 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_26 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_18_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_19_stat_bpd_mispredicted <= _T_28623 & _T_76 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_27 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_19_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_20_stat_bpd_mispredicted <= _T_28623 & _T_77 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_28 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_20_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_21_stat_bpd_mispredicted <= _T_28623 & _T_78 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_29 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_21_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_22_stat_bpd_mispredicted <= _T_28623 & _T_79 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_30 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_22_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_23_stat_bpd_mispredicted <= _T_28623 & _T_80 ? io_brinfo_bpd_mispredict : io_dis_valids_0 & _T_31 ?
                                io_dis_uops_0_stat_bpd_mispredicted : T_26182_23_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_26182_0_stat_bpd_made_pred <= _T_28623 & _T_57 ? io_brinfo_bpd_made_pred : ~io_dis_valids_0 | |rob_tail ?
                                T_26182_0_stat_bpd_made_pred : io_dis_uops_0_stat_bpd_made_pred;	// rob.scala:192:32, :347:34, :350:34, :406:72
    T_26182_1_stat_bpd_made_pred <= _T_28623 & _T_58 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_9 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_1_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_2_stat_bpd_made_pred <= _T_28623 & _T_59 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_10 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_2_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_3_stat_bpd_made_pred <= _T_28623 & _T_60 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_11 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_3_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_4_stat_bpd_made_pred <= _T_28623 & _T_61 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_12 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_4_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_5_stat_bpd_made_pred <= _T_28623 & _T_62 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_13 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_5_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_6_stat_bpd_made_pred <= _T_28623 & _T_63 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_14 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_6_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_7_stat_bpd_made_pred <= _T_28623 & _T_64 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_15 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_7_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_8_stat_bpd_made_pred <= _T_28623 & _T_65 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_16 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_8_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_9_stat_bpd_made_pred <= _T_28623 & _T_66 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_17 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_9_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_10_stat_bpd_made_pred <= _T_28623 & _T_67 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_18 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_10_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_11_stat_bpd_made_pred <= _T_28623 & _T_68 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_19 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_11_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_12_stat_bpd_made_pred <= _T_28623 & _T_69 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_20 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_12_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_13_stat_bpd_made_pred <= _T_28623 & _T_70 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_21 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_13_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_14_stat_bpd_made_pred <= _T_28623 & _T_71 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_22 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_14_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_15_stat_bpd_made_pred <= _T_28623 & _T_72 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_23 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_15_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_16_stat_bpd_made_pred <= _T_28623 & _T_73 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_24 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_16_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_17_stat_bpd_made_pred <= _T_28623 & _T_74 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_25 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_17_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_18_stat_bpd_made_pred <= _T_28623 & _T_75 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_26 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_18_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_19_stat_bpd_made_pred <= _T_28623 & _T_76 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_27 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_19_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_20_stat_bpd_made_pred <= _T_28623 & _T_77 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_28 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_20_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_21_stat_bpd_made_pred <= _T_28623 & _T_78 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_29 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_21_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_22_stat_bpd_made_pred <= _T_28623 & _T_79 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_30 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_22_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_23_stat_bpd_made_pred <= _T_28623 & _T_80 ? io_brinfo_bpd_made_pred : io_dis_valids_0 & _T_31 ?
                                io_dis_uops_0_stat_bpd_made_pred : T_26182_23_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_26182_0_br_mask <= ~_T_29370 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29368 ? T_26182_0_br_mask &
                                ~io_brinfo_mask : ~io_dis_valids_0 | |rob_tail ? T_26182_0_br_mask : io_dis_uops_0_br_mask;	// rob.scala:192:32, :347:34, :350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_1_br_mask <= ~_T_29472 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29470 ? T_26182_1_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_9 ? io_dis_uops_0_br_mask : T_26182_1_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_2_br_mask <= ~_T_29574 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29572 ? T_26182_2_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_10 ? io_dis_uops_0_br_mask : T_26182_2_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_3_br_mask <= ~_T_29676 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29674 ? T_26182_3_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_11 ? io_dis_uops_0_br_mask : T_26182_3_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_4_br_mask <= ~_T_29778 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29776 ? T_26182_4_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_12 ? io_dis_uops_0_br_mask : T_26182_4_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_5_br_mask <= ~_T_29880 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29878 ? T_26182_5_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_13 ? io_dis_uops_0_br_mask : T_26182_5_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_6_br_mask <= ~_T_29982 & io_brinfo_valid & ~io_brinfo_mispredict & _T_29980 ? T_26182_6_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_14 ? io_dis_uops_0_br_mask : T_26182_6_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_7_br_mask <= ~_T_30084 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30082 ? T_26182_7_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_15 ? io_dis_uops_0_br_mask : T_26182_7_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_8_br_mask <= ~_T_30186 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30184 ? T_26182_8_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_16 ? io_dis_uops_0_br_mask : T_26182_8_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_9_br_mask <= ~_T_30288 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30286 ? T_26182_9_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_17 ? io_dis_uops_0_br_mask : T_26182_9_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_10_br_mask <= ~_T_30390 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30388 ? T_26182_10_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_18 ? io_dis_uops_0_br_mask : T_26182_10_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_11_br_mask <= ~_T_30492 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30490 ? T_26182_11_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_19 ? io_dis_uops_0_br_mask : T_26182_11_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_12_br_mask <= ~_T_30594 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30592 ? T_26182_12_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_20 ? io_dis_uops_0_br_mask : T_26182_12_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_13_br_mask <= ~_T_30696 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30694 ? T_26182_13_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_21 ? io_dis_uops_0_br_mask : T_26182_13_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_14_br_mask <= ~_T_30798 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30796 ? T_26182_14_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_22 ? io_dis_uops_0_br_mask : T_26182_14_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_15_br_mask <= ~_T_30900 & io_brinfo_valid & ~io_brinfo_mispredict & _T_30898 ? T_26182_15_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_23 ? io_dis_uops_0_br_mask : T_26182_15_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_16_br_mask <= ~_T_31002 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31000 ? T_26182_16_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_24 ? io_dis_uops_0_br_mask : T_26182_16_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_17_br_mask <= ~_T_31104 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31102 ? T_26182_17_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_25 ? io_dis_uops_0_br_mask : T_26182_17_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_18_br_mask <= ~_T_31206 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31204 ? T_26182_18_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_26 ? io_dis_uops_0_br_mask : T_26182_18_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_19_br_mask <= ~_T_31308 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31306 ? T_26182_19_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_27 ? io_dis_uops_0_br_mask : T_26182_19_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_20_br_mask <= ~_T_31410 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31408 ? T_26182_20_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_28 ? io_dis_uops_0_br_mask : T_26182_20_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_21_br_mask <= ~_T_31512 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31510 ? T_26182_21_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_29 ? io_dis_uops_0_br_mask : T_26182_21_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_22_br_mask <= ~_T_31614 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31612 ? T_26182_22_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_30 ? io_dis_uops_0_br_mask : T_26182_22_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_23_br_mask <= ~_T_31716 & io_brinfo_valid & ~io_brinfo_mispredict & _T_31714 ? T_26182_23_br_mask &
                                ~io_brinfo_mask : io_dis_valids_0 & _T_31 ? io_dis_uops_0_br_mask : T_26182_23_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_26182_0_inst <= ~_T_32082 | |rob_tail ? (_T_3 ? (~(|rob_head) | _T_104 ? 32'h4033 : _T_32) : _T_104 ?
                                32'h4033 : _T_32) : 32'h4033;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :347:34, :357:33, :487:35, :500:28, :515:33, :519:33
    T_26182_1_inst <= _T_32082 & _T_9 ? 32'h4033 : _T_3 ? (_T_81 | _T_105 ? 32'h4033 : _T_33) : _T_105 ? 32'h4033
                                : _T_33;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_2_inst <= _T_32082 & _T_10 ? 32'h4033 : _T_3 ? (_T_82 | _T_106 ? 32'h4033 : _T_34) : _T_106 ?
                                32'h4033 : _T_34;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_3_inst <= _T_32082 & _T_11 ? 32'h4033 : _T_3 ? (_T_83 | _T_107 ? 32'h4033 : _T_35) : _T_107 ?
                                32'h4033 : _T_35;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_4_inst <= _T_32082 & _T_12 ? 32'h4033 : _T_3 ? (_T_84 | _T_108 ? 32'h4033 : _T_36) : _T_108 ?
                                32'h4033 : _T_36;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_5_inst <= _T_32082 & _T_13 ? 32'h4033 : _T_3 ? (_T_85 | _T_109 ? 32'h4033 : _T_37) : _T_109 ?
                                32'h4033 : _T_37;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_6_inst <= _T_32082 & _T_14 ? 32'h4033 : _T_3 ? (_T_86 | _T_110 ? 32'h4033 : _T_38) : _T_110 ?
                                32'h4033 : _T_38;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_7_inst <= _T_32082 & _T_15 ? 32'h4033 : _T_3 ? (_T_87 | _T_111 ? 32'h4033 : _T_39) : _T_111 ?
                                32'h4033 : _T_39;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_8_inst <= _T_32082 & _T_16 ? 32'h4033 : _T_3 ? (_T_88 | _T_112 ? 32'h4033 : _T_40) : _T_112 ?
                                32'h4033 : _T_40;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_9_inst <= _T_32082 & _T_17 ? 32'h4033 : _T_3 ? (_T_89 | _T_113 ? 32'h4033 : _T_41) : _T_113 ?
                                32'h4033 : _T_41;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_10_inst <= _T_32082 & _T_18 ? 32'h4033 : _T_3 ? (_T_90 | _T_114 ? 32'h4033 : _T_42) : _T_114 ?
                                32'h4033 : _T_42;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_11_inst <= _T_32082 & _T_19 ? 32'h4033 : _T_3 ? (_T_91 | _T_115 ? 32'h4033 : _T_43) : _T_115 ?
                                32'h4033 : _T_43;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_12_inst <= _T_32082 & _T_20 ? 32'h4033 : _T_3 ? (_T_92 | _T_116 ? 32'h4033 : _T_44) : _T_116 ?
                                32'h4033 : _T_44;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_13_inst <= _T_32082 & _T_21 ? 32'h4033 : _T_3 ? (_T_93 | _T_117 ? 32'h4033 : _T_45) : _T_117 ?
                                32'h4033 : _T_45;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_14_inst <= _T_32082 & _T_22 ? 32'h4033 : _T_3 ? (_T_94 | _T_118 ? 32'h4033 : _T_46) : _T_118 ?
                                32'h4033 : _T_46;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_15_inst <= _T_32082 & _T_23 ? 32'h4033 : _T_3 ? (_T_95 | _T_119 ? 32'h4033 : _T_47) : _T_119 ?
                                32'h4033 : _T_47;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_16_inst <= _T_32082 & _T_24 ? 32'h4033 : _T_3 ? (_T_96 | _T_120 ? 32'h4033 : _T_48) : _T_120 ?
                                32'h4033 : _T_48;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_17_inst <= _T_32082 & _T_25 ? 32'h4033 : _T_3 ? (_T_97 | _T_121 ? 32'h4033 : _T_49) : _T_121 ?
                                32'h4033 : _T_49;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_18_inst <= _T_32082 & _T_26 ? 32'h4033 : _T_3 ? (_T_98 | _T_122 ? 32'h4033 : _T_50) : _T_122 ?
                                32'h4033 : _T_50;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_19_inst <= _T_32082 & _T_27 ? 32'h4033 : _T_3 ? (_T_99 | _T_123 ? 32'h4033 : _T_51) : _T_123 ?
                                32'h4033 : _T_51;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_20_inst <= _T_32082 & _T_28 ? 32'h4033 : _T_3 ? (_T_100 | _T_124 ? 32'h4033 : _T_52) : _T_124 ?
                                32'h4033 : _T_52;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_21_inst <= _T_32082 & _T_29 ? 32'h4033 : _T_3 ? (_T_101 | _T_125 ? 32'h4033 : _T_53) : _T_125 ?
                                32'h4033 : _T_53;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_22_inst <= _T_32082 & _T_30 ? 32'h4033 : _T_3 ? (_T_102 | _T_126 ? 32'h4033 : _T_54) : _T_126 ?
                                32'h4033 : _T_54;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_26182_23_inst <= _T_32082 & _T_31 ? 32'h4033 : _T_3 ? (_T_103 | _T_127 ? 32'h4033 : _T_55) : _T_127 ?
                                32'h4033 : _T_55;	// rob.scala:357:33, :487:35, :515:33, :519:33
    `ifndef SYNTHESIS	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_32357)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_32357)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_32369)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_32369)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
      if (`PRINTF_COND_ & ~_T_32561)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_32561)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_32573)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_32573)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
    `endif
    T_26182_0_debug_wdata <= _T_32579 & _T_176 ? io_debug_wb_wdata_2 : _T_32375 & _T_152 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_128 ? io_debug_wb_wdata_0 : ~io_dis_valids_0 | |rob_tail ?
                                T_26182_0_debug_wdata : io_dis_uops_0_debug_wdata;	// rob.scala:192:32, :347:34, :350:34, :531:53
    T_26182_1_debug_wdata <= _T_32579 & _T_177 ? io_debug_wb_wdata_2 : _T_32375 & _T_153 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_129 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_9 ?
                                io_dis_uops_0_debug_wdata : T_26182_1_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_2_debug_wdata <= _T_32579 & _T_178 ? io_debug_wb_wdata_2 : _T_32375 & _T_154 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_130 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_10 ?
                                io_dis_uops_0_debug_wdata : T_26182_2_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_3_debug_wdata <= _T_32579 & _T_179 ? io_debug_wb_wdata_2 : _T_32375 & _T_155 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_131 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_11 ?
                                io_dis_uops_0_debug_wdata : T_26182_3_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_4_debug_wdata <= _T_32579 & _T_180 ? io_debug_wb_wdata_2 : _T_32375 & _T_156 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_132 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_12 ?
                                io_dis_uops_0_debug_wdata : T_26182_4_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_5_debug_wdata <= _T_32579 & _T_181 ? io_debug_wb_wdata_2 : _T_32375 & _T_157 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_133 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_13 ?
                                io_dis_uops_0_debug_wdata : T_26182_5_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_6_debug_wdata <= _T_32579 & _T_182 ? io_debug_wb_wdata_2 : _T_32375 & _T_158 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_134 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_14 ?
                                io_dis_uops_0_debug_wdata : T_26182_6_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_7_debug_wdata <= _T_32579 & _T_183 ? io_debug_wb_wdata_2 : _T_32375 & _T_159 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_135 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_15 ?
                                io_dis_uops_0_debug_wdata : T_26182_7_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_8_debug_wdata <= _T_32579 & _T_184 ? io_debug_wb_wdata_2 : _T_32375 & _T_160 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_136 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_16 ?
                                io_dis_uops_0_debug_wdata : T_26182_8_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_9_debug_wdata <= _T_32579 & _T_185 ? io_debug_wb_wdata_2 : _T_32375 & _T_161 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_137 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_17 ?
                                io_dis_uops_0_debug_wdata : T_26182_9_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_10_debug_wdata <= _T_32579 & _T_186 ? io_debug_wb_wdata_2 : _T_32375 & _T_162 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_138 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_18 ?
                                io_dis_uops_0_debug_wdata : T_26182_10_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_11_debug_wdata <= _T_32579 & _T_187 ? io_debug_wb_wdata_2 : _T_32375 & _T_163 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_139 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_19 ?
                                io_dis_uops_0_debug_wdata : T_26182_11_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_12_debug_wdata <= _T_32579 & _T_188 ? io_debug_wb_wdata_2 : _T_32375 & _T_164 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_140 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_20 ?
                                io_dis_uops_0_debug_wdata : T_26182_12_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_13_debug_wdata <= _T_32579 & _T_189 ? io_debug_wb_wdata_2 : _T_32375 & _T_165 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_141 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_21 ?
                                io_dis_uops_0_debug_wdata : T_26182_13_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_14_debug_wdata <= _T_32579 & _T_190 ? io_debug_wb_wdata_2 : _T_32375 & _T_166 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_142 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_22 ?
                                io_dis_uops_0_debug_wdata : T_26182_14_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_15_debug_wdata <= _T_32579 & _T_191 ? io_debug_wb_wdata_2 : _T_32375 & _T_167 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_143 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_23 ?
                                io_dis_uops_0_debug_wdata : T_26182_15_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_16_debug_wdata <= _T_32579 & _T_192 ? io_debug_wb_wdata_2 : _T_32375 & _T_168 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_144 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_24 ?
                                io_dis_uops_0_debug_wdata : T_26182_16_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_17_debug_wdata <= _T_32579 & _T_193 ? io_debug_wb_wdata_2 : _T_32375 & _T_169 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_145 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_25 ?
                                io_dis_uops_0_debug_wdata : T_26182_17_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_18_debug_wdata <= _T_32579 & _T_194 ? io_debug_wb_wdata_2 : _T_32375 & _T_170 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_146 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_26 ?
                                io_dis_uops_0_debug_wdata : T_26182_18_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_19_debug_wdata <= _T_32579 & _T_195 ? io_debug_wb_wdata_2 : _T_32375 & _T_171 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_147 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_27 ?
                                io_dis_uops_0_debug_wdata : T_26182_19_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_20_debug_wdata <= _T_32579 & _T_196 ? io_debug_wb_wdata_2 : _T_32375 & _T_172 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_148 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_28 ?
                                io_dis_uops_0_debug_wdata : T_26182_20_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_21_debug_wdata <= _T_32579 & _T_197 ? io_debug_wb_wdata_2 : _T_32375 & _T_173 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_149 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_29 ?
                                io_dis_uops_0_debug_wdata : T_26182_21_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_22_debug_wdata <= _T_32579 & _T_198 ? io_debug_wb_wdata_2 : _T_32375 & _T_174 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_150 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_30 ?
                                io_dis_uops_0_debug_wdata : T_26182_22_debug_wdata;	// rob.scala:350:34, :531:53
    T_26182_23_debug_wdata <= _T_32579 & _T_199 ? io_debug_wb_wdata_2 : _T_32375 & _T_175 ? io_debug_wb_wdata_1 :
                                _T_32171 & _T_151 ? io_debug_wb_wdata_0 : io_dis_valids_0 & _T_31 ?
                                io_dis_uops_0_debug_wdata : T_26182_23_debug_wdata;	// rob.scala:350:34, :531:53
    `ifndef SYNTHESIS	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_32765)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_32765)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_32777)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_32777)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
    `endif
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (~(~io_dis_valids_1 | |rob_tail))	// rob.scala:192:32, :347:34, :350:34
      T_38110_0_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_9)	// rob.scala:350:34
      T_38110_1_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_10)	// rob.scala:350:34
      T_38110_2_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_11)	// rob.scala:350:34
      T_38110_3_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_12)	// rob.scala:350:34
      T_38110_4_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_13)	// rob.scala:350:34
      T_38110_5_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_14)	// rob.scala:350:34
      T_38110_6_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_15)	// rob.scala:350:34
      T_38110_7_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_16)	// rob.scala:350:34
      T_38110_8_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_17)	// rob.scala:350:34
      T_38110_9_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_18)	// rob.scala:350:34
      T_38110_10_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_19)	// rob.scala:350:34
      T_38110_11_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_20)	// rob.scala:350:34
      T_38110_12_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_21)	// rob.scala:350:34
      T_38110_13_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_22)	// rob.scala:350:34
      T_38110_14_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_23)	// rob.scala:350:34
      T_38110_15_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_24)	// rob.scala:350:34
      T_38110_16_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_25)	// rob.scala:350:34
      T_38110_17_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_26)	// rob.scala:350:34
      T_38110_18_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_27)	// rob.scala:350:34
      T_38110_19_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_28)	// rob.scala:350:34
      T_38110_20_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_29)	// rob.scala:350:34
      T_38110_21_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_30)	// rob.scala:350:34
      T_38110_22_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_valid <= io_dis_uops_1_valid;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_iw_state <= io_dis_uops_1_iw_state;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_uopc <= io_dis_uops_1_uopc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_pc <= io_dis_uops_1_pc;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_fu_code <= io_dis_uops_1_fu_code;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_br_type <= io_dis_uops_1_ctrl_br_type;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_op1_sel <= io_dis_uops_1_ctrl_op1_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_op2_sel <= io_dis_uops_1_ctrl_op2_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_imm_sel <= io_dis_uops_1_ctrl_imm_sel;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_op_fcn <= io_dis_uops_1_ctrl_op_fcn;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_fcn_dw <= io_dis_uops_1_ctrl_fcn_dw;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_rf_wen <= io_dis_uops_1_ctrl_rf_wen;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_csr_cmd <= io_dis_uops_1_ctrl_csr_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_is_load <= io_dis_uops_1_ctrl_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_is_sta <= io_dis_uops_1_ctrl_is_sta;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ctrl_is_std <= io_dis_uops_1_ctrl_is_std;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_wakeup_delay <= io_dis_uops_1_wakeup_delay;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_allocate_brtag <= io_dis_uops_1_allocate_brtag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_br_or_jmp <= io_dis_uops_1_is_br_or_jmp;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_jump <= io_dis_uops_1_is_jump;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_jal <= io_dis_uops_1_is_jal;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_ret <= io_dis_uops_1_is_ret;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_call <= io_dis_uops_1_is_call;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_tag <= io_dis_uops_1_br_tag;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_prediction_bpd_predict_val <= io_dis_uops_1_br_prediction_bpd_predict_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_prediction_bpd_predict_taken <= io_dis_uops_1_br_prediction_bpd_predict_taken;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_prediction_btb_hit <= io_dis_uops_1_br_prediction_btb_hit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_prediction_btb_predicted <= io_dis_uops_1_br_prediction_btb_predicted;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_br_prediction_is_br_or_jalr <= io_dis_uops_1_br_prediction_is_br_or_jalr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_fetch_pc_lob <= io_dis_uops_1_fetch_pc_lob;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_imm_packed <= io_dis_uops_1_imm_packed;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_csr_addr <= io_dis_uops_1_csr_addr;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_rob_idx <= io_dis_uops_1_rob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ldq_idx <= io_dis_uops_1_ldq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_stq_idx <= io_dis_uops_1_stq_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_brob_idx <= io_dis_uops_1_brob_idx;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_pdst <= io_dis_uops_1_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_pop1 <= io_dis_uops_1_pop1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_pop2 <= io_dis_uops_1_pop2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_pop3 <= io_dis_uops_1_pop3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_prs1_busy <= io_dis_uops_1_prs1_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_prs2_busy <= io_dis_uops_1_prs2_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_prs3_busy <= io_dis_uops_1_prs3_busy;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_stale_pdst <= io_dis_uops_1_stale_pdst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_exception <= io_dis_uops_1_exception;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_exc_cause <= io_dis_uops_1_exc_cause;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_bypassable <= io_dis_uops_1_bypassable;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_mem_cmd <= io_dis_uops_1_mem_cmd;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_mem_typ <= io_dis_uops_1_mem_typ;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_fence <= io_dis_uops_1_is_fence;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_fencei <= io_dis_uops_1_is_fencei;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_store <= io_dis_uops_1_is_store;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_amo <= io_dis_uops_1_is_amo;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_load <= io_dis_uops_1_is_load;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_is_unique <= io_dis_uops_1_is_unique;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_flush_on_commit <= io_dis_uops_1_flush_on_commit;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ldst <= io_dis_uops_1_ldst;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_lrs1 <= io_dis_uops_1_lrs1;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_lrs2 <= io_dis_uops_1_lrs2;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_lrs3 <= io_dis_uops_1_lrs3;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_ldst_val <= io_dis_uops_1_ldst_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_dst_rtype <= io_dis_uops_1_dst_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_lrs1_rtype <= io_dis_uops_1_lrs1_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_lrs2_rtype <= io_dis_uops_1_lrs2_rtype;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_frs3_en <= io_dis_uops_1_frs3_en;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_fp_val <= io_dis_uops_1_fp_val;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_fp_single <= io_dis_uops_1_fp_single;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_xcpt_if <= io_dis_uops_1_xcpt_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_replay_if <= io_dis_uops_1_replay_if;	// rob.scala:350:34
    if (io_dis_valids_1 & _T_31)	// rob.scala:350:34
      T_38110_23_debug_events_fetch_seq <= io_dis_uops_1_debug_events_fetch_seq;	// rob.scala:350:34
    T_38110_0_stat_brjmp_mispredicted <= _T_40551 & _T_57 ? io_brinfo_mispredict : io_dis_valids_1 ? |rob_tail & (|rob_tail ?
                                T_38110_0_stat_brjmp_mispredicted : io_dis_uops_1_stat_brjmp_mispredicted) :
                                T_38110_0_stat_brjmp_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :353:52, :402:72
    T_38110_1_stat_brjmp_mispredicted <= _T_40551 & _T_58 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_9 & (_T_9 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_1_stat_brjmp_mispredicted) :
                                T_38110_1_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_2_stat_brjmp_mispredicted <= _T_40551 & _T_59 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_10 & (_T_10 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_2_stat_brjmp_mispredicted) :
                                T_38110_2_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_3_stat_brjmp_mispredicted <= _T_40551 & _T_60 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_11 & (_T_11 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_3_stat_brjmp_mispredicted) :
                                T_38110_3_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_4_stat_brjmp_mispredicted <= _T_40551 & _T_61 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_12 & (_T_12 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_4_stat_brjmp_mispredicted) :
                                T_38110_4_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_5_stat_brjmp_mispredicted <= _T_40551 & _T_62 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_13 & (_T_13 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_5_stat_brjmp_mispredicted) :
                                T_38110_5_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_6_stat_brjmp_mispredicted <= _T_40551 & _T_63 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_14 & (_T_14 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_6_stat_brjmp_mispredicted) :
                                T_38110_6_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_7_stat_brjmp_mispredicted <= _T_40551 & _T_64 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_15 & (_T_15 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_7_stat_brjmp_mispredicted) :
                                T_38110_7_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_8_stat_brjmp_mispredicted <= _T_40551 & _T_65 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_16 & (_T_16 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_8_stat_brjmp_mispredicted) :
                                T_38110_8_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_9_stat_brjmp_mispredicted <= _T_40551 & _T_66 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_17 & (_T_17 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_9_stat_brjmp_mispredicted) :
                                T_38110_9_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_10_stat_brjmp_mispredicted <= _T_40551 & _T_67 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_18 & (_T_18 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_10_stat_brjmp_mispredicted) :
                                T_38110_10_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_11_stat_brjmp_mispredicted <= _T_40551 & _T_68 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_19 & (_T_19 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_11_stat_brjmp_mispredicted) :
                                T_38110_11_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_12_stat_brjmp_mispredicted <= _T_40551 & _T_69 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_20 & (_T_20 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_12_stat_brjmp_mispredicted) :
                                T_38110_12_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_13_stat_brjmp_mispredicted <= _T_40551 & _T_70 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_21 & (_T_21 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_13_stat_brjmp_mispredicted) :
                                T_38110_13_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_14_stat_brjmp_mispredicted <= _T_40551 & _T_71 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_22 & (_T_22 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_14_stat_brjmp_mispredicted) :
                                T_38110_14_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_15_stat_brjmp_mispredicted <= _T_40551 & _T_72 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_23 & (_T_23 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_15_stat_brjmp_mispredicted) :
                                T_38110_15_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_16_stat_brjmp_mispredicted <= _T_40551 & _T_73 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_24 & (_T_24 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_16_stat_brjmp_mispredicted) :
                                T_38110_16_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_17_stat_brjmp_mispredicted <= _T_40551 & _T_74 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_25 & (_T_25 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_17_stat_brjmp_mispredicted) :
                                T_38110_17_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_18_stat_brjmp_mispredicted <= _T_40551 & _T_75 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_26 & (_T_26 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_18_stat_brjmp_mispredicted) :
                                T_38110_18_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_19_stat_brjmp_mispredicted <= _T_40551 & _T_76 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_27 & (_T_27 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_19_stat_brjmp_mispredicted) :
                                T_38110_19_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_20_stat_brjmp_mispredicted <= _T_40551 & _T_77 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_28 & (_T_28 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_20_stat_brjmp_mispredicted) :
                                T_38110_20_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_21_stat_brjmp_mispredicted <= _T_40551 & _T_78 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_29 & (_T_29 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_21_stat_brjmp_mispredicted) :
                                T_38110_21_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_22_stat_brjmp_mispredicted <= _T_40551 & _T_79 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_30 & (_T_30 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_22_stat_brjmp_mispredicted) :
                                T_38110_22_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_23_stat_brjmp_mispredicted <= _T_40551 & _T_80 ? io_brinfo_mispredict : io_dis_valids_1 ? ~_T_31 & (_T_31 ?
                                io_dis_uops_1_stat_brjmp_mispredicted : T_38110_23_stat_brjmp_mispredicted) :
                                T_38110_23_stat_brjmp_mispredicted;	// rob.scala:350:34, :353:52, :402:72
    T_38110_0_stat_btb_mispredicted <= _T_40551 & _T_57 ? io_brinfo_btb_mispredict : ~io_dis_valids_1 | |rob_tail ?
                                T_38110_0_stat_btb_mispredicted : io_dis_uops_1_stat_btb_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :403:72
    T_38110_1_stat_btb_mispredicted <= _T_40551 & _T_58 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_9 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_1_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_2_stat_btb_mispredicted <= _T_40551 & _T_59 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_10 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_2_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_3_stat_btb_mispredicted <= _T_40551 & _T_60 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_11 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_3_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_4_stat_btb_mispredicted <= _T_40551 & _T_61 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_12 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_4_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_5_stat_btb_mispredicted <= _T_40551 & _T_62 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_13 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_5_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_6_stat_btb_mispredicted <= _T_40551 & _T_63 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_14 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_6_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_7_stat_btb_mispredicted <= _T_40551 & _T_64 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_15 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_7_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_8_stat_btb_mispredicted <= _T_40551 & _T_65 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_16 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_8_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_9_stat_btb_mispredicted <= _T_40551 & _T_66 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_17 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_9_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_10_stat_btb_mispredicted <= _T_40551 & _T_67 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_18 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_10_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_11_stat_btb_mispredicted <= _T_40551 & _T_68 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_19 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_11_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_12_stat_btb_mispredicted <= _T_40551 & _T_69 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_20 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_12_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_13_stat_btb_mispredicted <= _T_40551 & _T_70 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_21 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_13_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_14_stat_btb_mispredicted <= _T_40551 & _T_71 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_22 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_14_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_15_stat_btb_mispredicted <= _T_40551 & _T_72 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_23 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_15_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_16_stat_btb_mispredicted <= _T_40551 & _T_73 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_24 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_16_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_17_stat_btb_mispredicted <= _T_40551 & _T_74 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_25 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_17_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_18_stat_btb_mispredicted <= _T_40551 & _T_75 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_26 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_18_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_19_stat_btb_mispredicted <= _T_40551 & _T_76 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_27 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_19_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_20_stat_btb_mispredicted <= _T_40551 & _T_77 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_28 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_20_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_21_stat_btb_mispredicted <= _T_40551 & _T_78 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_29 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_21_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_22_stat_btb_mispredicted <= _T_40551 & _T_79 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_30 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_22_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_23_stat_btb_mispredicted <= _T_40551 & _T_80 ? io_brinfo_btb_mispredict : io_dis_valids_1 & _T_31 ?
                                io_dis_uops_1_stat_btb_mispredicted : T_38110_23_stat_btb_mispredicted;	// rob.scala:350:34, :403:72
    T_38110_0_stat_btb_made_pred <= _T_40551 & _T_57 ? io_brinfo_btb_made_pred : ~io_dis_valids_1 | |rob_tail ?
                                T_38110_0_stat_btb_made_pred : io_dis_uops_1_stat_btb_made_pred;	// rob.scala:192:32, :347:34, :350:34, :404:72
    T_38110_1_stat_btb_made_pred <= _T_40551 & _T_58 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_9 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_1_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_2_stat_btb_made_pred <= _T_40551 & _T_59 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_10 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_2_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_3_stat_btb_made_pred <= _T_40551 & _T_60 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_11 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_3_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_4_stat_btb_made_pred <= _T_40551 & _T_61 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_12 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_4_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_5_stat_btb_made_pred <= _T_40551 & _T_62 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_13 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_5_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_6_stat_btb_made_pred <= _T_40551 & _T_63 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_14 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_6_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_7_stat_btb_made_pred <= _T_40551 & _T_64 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_15 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_7_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_8_stat_btb_made_pred <= _T_40551 & _T_65 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_16 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_8_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_9_stat_btb_made_pred <= _T_40551 & _T_66 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_17 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_9_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_10_stat_btb_made_pred <= _T_40551 & _T_67 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_18 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_10_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_11_stat_btb_made_pred <= _T_40551 & _T_68 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_19 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_11_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_12_stat_btb_made_pred <= _T_40551 & _T_69 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_20 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_12_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_13_stat_btb_made_pred <= _T_40551 & _T_70 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_21 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_13_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_14_stat_btb_made_pred <= _T_40551 & _T_71 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_22 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_14_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_15_stat_btb_made_pred <= _T_40551 & _T_72 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_23 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_15_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_16_stat_btb_made_pred <= _T_40551 & _T_73 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_24 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_16_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_17_stat_btb_made_pred <= _T_40551 & _T_74 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_25 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_17_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_18_stat_btb_made_pred <= _T_40551 & _T_75 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_26 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_18_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_19_stat_btb_made_pred <= _T_40551 & _T_76 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_27 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_19_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_20_stat_btb_made_pred <= _T_40551 & _T_77 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_28 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_20_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_21_stat_btb_made_pred <= _T_40551 & _T_78 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_29 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_21_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_22_stat_btb_made_pred <= _T_40551 & _T_79 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_30 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_22_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_23_stat_btb_made_pred <= _T_40551 & _T_80 ? io_brinfo_btb_made_pred : io_dis_valids_1 & _T_31 ?
                                io_dis_uops_1_stat_btb_made_pred : T_38110_23_stat_btb_made_pred;	// rob.scala:350:34, :404:72
    T_38110_0_stat_bpd_mispredicted <= _T_40551 & _T_57 ? io_brinfo_bpd_mispredict : ~io_dis_valids_1 | |rob_tail ?
                                T_38110_0_stat_bpd_mispredicted : io_dis_uops_1_stat_bpd_mispredicted;	// rob.scala:192:32, :347:34, :350:34, :405:72
    T_38110_1_stat_bpd_mispredicted <= _T_40551 & _T_58 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_9 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_1_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_2_stat_bpd_mispredicted <= _T_40551 & _T_59 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_10 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_2_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_3_stat_bpd_mispredicted <= _T_40551 & _T_60 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_11 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_3_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_4_stat_bpd_mispredicted <= _T_40551 & _T_61 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_12 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_4_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_5_stat_bpd_mispredicted <= _T_40551 & _T_62 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_13 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_5_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_6_stat_bpd_mispredicted <= _T_40551 & _T_63 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_14 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_6_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_7_stat_bpd_mispredicted <= _T_40551 & _T_64 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_15 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_7_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_8_stat_bpd_mispredicted <= _T_40551 & _T_65 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_16 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_8_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_9_stat_bpd_mispredicted <= _T_40551 & _T_66 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_17 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_9_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_10_stat_bpd_mispredicted <= _T_40551 & _T_67 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_18 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_10_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_11_stat_bpd_mispredicted <= _T_40551 & _T_68 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_19 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_11_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_12_stat_bpd_mispredicted <= _T_40551 & _T_69 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_20 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_12_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_13_stat_bpd_mispredicted <= _T_40551 & _T_70 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_21 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_13_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_14_stat_bpd_mispredicted <= _T_40551 & _T_71 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_22 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_14_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_15_stat_bpd_mispredicted <= _T_40551 & _T_72 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_23 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_15_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_16_stat_bpd_mispredicted <= _T_40551 & _T_73 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_24 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_16_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_17_stat_bpd_mispredicted <= _T_40551 & _T_74 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_25 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_17_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_18_stat_bpd_mispredicted <= _T_40551 & _T_75 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_26 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_18_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_19_stat_bpd_mispredicted <= _T_40551 & _T_76 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_27 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_19_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_20_stat_bpd_mispredicted <= _T_40551 & _T_77 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_28 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_20_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_21_stat_bpd_mispredicted <= _T_40551 & _T_78 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_29 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_21_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_22_stat_bpd_mispredicted <= _T_40551 & _T_79 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_30 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_22_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_23_stat_bpd_mispredicted <= _T_40551 & _T_80 ? io_brinfo_bpd_mispredict : io_dis_valids_1 & _T_31 ?
                                io_dis_uops_1_stat_bpd_mispredicted : T_38110_23_stat_bpd_mispredicted;	// rob.scala:350:34, :405:72
    T_38110_0_stat_bpd_made_pred <= _T_40551 & _T_57 ? io_brinfo_bpd_made_pred : ~io_dis_valids_1 | |rob_tail ?
                                T_38110_0_stat_bpd_made_pred : io_dis_uops_1_stat_bpd_made_pred;	// rob.scala:192:32, :347:34, :350:34, :406:72
    T_38110_1_stat_bpd_made_pred <= _T_40551 & _T_58 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_9 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_1_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_2_stat_bpd_made_pred <= _T_40551 & _T_59 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_10 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_2_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_3_stat_bpd_made_pred <= _T_40551 & _T_60 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_11 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_3_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_4_stat_bpd_made_pred <= _T_40551 & _T_61 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_12 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_4_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_5_stat_bpd_made_pred <= _T_40551 & _T_62 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_13 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_5_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_6_stat_bpd_made_pred <= _T_40551 & _T_63 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_14 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_6_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_7_stat_bpd_made_pred <= _T_40551 & _T_64 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_15 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_7_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_8_stat_bpd_made_pred <= _T_40551 & _T_65 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_16 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_8_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_9_stat_bpd_made_pred <= _T_40551 & _T_66 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_17 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_9_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_10_stat_bpd_made_pred <= _T_40551 & _T_67 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_18 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_10_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_11_stat_bpd_made_pred <= _T_40551 & _T_68 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_19 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_11_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_12_stat_bpd_made_pred <= _T_40551 & _T_69 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_20 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_12_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_13_stat_bpd_made_pred <= _T_40551 & _T_70 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_21 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_13_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_14_stat_bpd_made_pred <= _T_40551 & _T_71 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_22 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_14_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_15_stat_bpd_made_pred <= _T_40551 & _T_72 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_23 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_15_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_16_stat_bpd_made_pred <= _T_40551 & _T_73 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_24 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_16_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_17_stat_bpd_made_pred <= _T_40551 & _T_74 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_25 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_17_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_18_stat_bpd_made_pred <= _T_40551 & _T_75 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_26 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_18_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_19_stat_bpd_made_pred <= _T_40551 & _T_76 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_27 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_19_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_20_stat_bpd_made_pred <= _T_40551 & _T_77 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_28 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_20_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_21_stat_bpd_made_pred <= _T_40551 & _T_78 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_29 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_21_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_22_stat_bpd_made_pred <= _T_40551 & _T_79 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_30 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_22_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_23_stat_bpd_made_pred <= _T_40551 & _T_80 ? io_brinfo_bpd_made_pred : io_dis_valids_1 & _T_31 ?
                                io_dis_uops_1_stat_bpd_made_pred : T_38110_23_stat_bpd_made_pred;	// rob.scala:350:34, :406:72
    T_38110_0_br_mask <= ~_T_41298 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41296 ? T_38110_0_br_mask &
                                ~io_brinfo_mask : ~io_dis_valids_1 | |rob_tail ? T_38110_0_br_mask : io_dis_uops_1_br_mask;	// rob.scala:192:32, :347:34, :350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_1_br_mask <= ~_T_41400 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41398 ? T_38110_1_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_9 ? io_dis_uops_1_br_mask : T_38110_1_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_2_br_mask <= ~_T_41502 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41500 ? T_38110_2_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_10 ? io_dis_uops_1_br_mask : T_38110_2_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_3_br_mask <= ~_T_41604 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41602 ? T_38110_3_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_11 ? io_dis_uops_1_br_mask : T_38110_3_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_4_br_mask <= ~_T_41706 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41704 ? T_38110_4_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_12 ? io_dis_uops_1_br_mask : T_38110_4_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_5_br_mask <= ~_T_41808 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41806 ? T_38110_5_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_13 ? io_dis_uops_1_br_mask : T_38110_5_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_6_br_mask <= ~_T_41910 & io_brinfo_valid & ~io_brinfo_mispredict & _T_41908 ? T_38110_6_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_14 ? io_dis_uops_1_br_mask : T_38110_6_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_7_br_mask <= ~_T_42012 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42010 ? T_38110_7_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_15 ? io_dis_uops_1_br_mask : T_38110_7_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_8_br_mask <= ~_T_42114 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42112 ? T_38110_8_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_16 ? io_dis_uops_1_br_mask : T_38110_8_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_9_br_mask <= ~_T_42216 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42214 ? T_38110_9_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_17 ? io_dis_uops_1_br_mask : T_38110_9_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_10_br_mask <= ~_T_42318 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42316 ? T_38110_10_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_18 ? io_dis_uops_1_br_mask : T_38110_10_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_11_br_mask <= ~_T_42420 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42418 ? T_38110_11_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_19 ? io_dis_uops_1_br_mask : T_38110_11_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_12_br_mask <= ~_T_42522 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42520 ? T_38110_12_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_20 ? io_dis_uops_1_br_mask : T_38110_12_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_13_br_mask <= ~_T_42624 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42622 ? T_38110_13_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_21 ? io_dis_uops_1_br_mask : T_38110_13_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_14_br_mask <= ~_T_42726 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42724 ? T_38110_14_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_22 ? io_dis_uops_1_br_mask : T_38110_14_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_15_br_mask <= ~_T_42828 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42826 ? T_38110_15_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_23 ? io_dis_uops_1_br_mask : T_38110_15_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_16_br_mask <= ~_T_42930 & io_brinfo_valid & ~io_brinfo_mispredict & _T_42928 ? T_38110_16_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_24 ? io_dis_uops_1_br_mask : T_38110_16_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_17_br_mask <= ~_T_43032 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43030 ? T_38110_17_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_25 ? io_dis_uops_1_br_mask : T_38110_17_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_18_br_mask <= ~_T_43134 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43132 ? T_38110_18_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_26 ? io_dis_uops_1_br_mask : T_38110_18_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_19_br_mask <= ~_T_43236 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43234 ? T_38110_19_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_27 ? io_dis_uops_1_br_mask : T_38110_19_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_20_br_mask <= ~_T_43338 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43336 ? T_38110_20_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_28 ? io_dis_uops_1_br_mask : T_38110_20_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_21_br_mask <= ~_T_43440 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43438 ? T_38110_21_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_29 ? io_dis_uops_1_br_mask : T_38110_21_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_22_br_mask <= ~_T_43542 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43540 ? T_38110_22_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_30 ? io_dis_uops_1_br_mask : T_38110_22_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_23_br_mask <= ~_T_43644 & io_brinfo_valid & ~io_brinfo_mispredict & _T_43642 ? T_38110_23_br_mask &
                                ~io_brinfo_mask : io_dis_valids_1 & _T_31 ? io_dis_uops_1_br_mask : T_38110_23_br_mask;	// rob.scala:350:34, :485:10, :489:40, :490:10, :492:{32,44,46}
    T_38110_0_inst <= ~_T_44010 | |rob_tail ? (_T_4 ? (~(|rob_head) | _T_225 ? 32'h4033 : _T_200) : _T_225 ?
                                32'h4033 : _T_200) : 32'h4033;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :347:34, :357:33, :487:35, :500:28, :515:33, :519:33
    T_38110_1_inst <= _T_44010 & _T_9 ? 32'h4033 : _T_4 ? (_T_81 | _T_226 ? 32'h4033 : _T_201) : _T_226 ?
                                32'h4033 : _T_201;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_2_inst <= _T_44010 & _T_10 ? 32'h4033 : _T_4 ? (_T_82 | _T_227 ? 32'h4033 : _T_202) : _T_227 ?
                                32'h4033 : _T_202;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_3_inst <= _T_44010 & _T_11 ? 32'h4033 : _T_4 ? (_T_83 | _T_228 ? 32'h4033 : _T_203) : _T_228 ?
                                32'h4033 : _T_203;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_4_inst <= _T_44010 & _T_12 ? 32'h4033 : _T_4 ? (_T_84 | _T_229 ? 32'h4033 : _T_204) : _T_229 ?
                                32'h4033 : _T_204;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_5_inst <= _T_44010 & _T_13 ? 32'h4033 : _T_4 ? (_T_85 | _T_230 ? 32'h4033 : _T_205) : _T_230 ?
                                32'h4033 : _T_205;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_6_inst <= _T_44010 & _T_14 ? 32'h4033 : _T_4 ? (_T_86 | _T_231 ? 32'h4033 : _T_206) : _T_231 ?
                                32'h4033 : _T_206;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_7_inst <= _T_44010 & _T_15 ? 32'h4033 : _T_4 ? (_T_87 | _T_232 ? 32'h4033 : _T_207) : _T_232 ?
                                32'h4033 : _T_207;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_8_inst <= _T_44010 & _T_16 ? 32'h4033 : _T_4 ? (_T_88 | _T_233 ? 32'h4033 : _T_208) : _T_233 ?
                                32'h4033 : _T_208;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_9_inst <= _T_44010 & _T_17 ? 32'h4033 : _T_4 ? (_T_89 | _T_234 ? 32'h4033 : _T_209) : _T_234 ?
                                32'h4033 : _T_209;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_10_inst <= _T_44010 & _T_18 ? 32'h4033 : _T_4 ? (_T_90 | _T_235 ? 32'h4033 : _T_210) : _T_235 ?
                                32'h4033 : _T_210;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_11_inst <= _T_44010 & _T_19 ? 32'h4033 : _T_4 ? (_T_91 | _T_236 ? 32'h4033 : _T_211) : _T_236 ?
                                32'h4033 : _T_211;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_12_inst <= _T_44010 & _T_20 ? 32'h4033 : _T_4 ? (_T_92 | _T_237 ? 32'h4033 : _T_212) : _T_237 ?
                                32'h4033 : _T_212;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_13_inst <= _T_44010 & _T_21 ? 32'h4033 : _T_4 ? (_T_93 | _T_238 ? 32'h4033 : _T_213) : _T_238 ?
                                32'h4033 : _T_213;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_14_inst <= _T_44010 & _T_22 ? 32'h4033 : _T_4 ? (_T_94 | _T_239 ? 32'h4033 : _T_214) : _T_239 ?
                                32'h4033 : _T_214;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_15_inst <= _T_44010 & _T_23 ? 32'h4033 : _T_4 ? (_T_95 | _T_240 ? 32'h4033 : _T_215) : _T_240 ?
                                32'h4033 : _T_215;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_16_inst <= _T_44010 & _T_24 ? 32'h4033 : _T_4 ? (_T_96 | _T_241 ? 32'h4033 : _T_216) : _T_241 ?
                                32'h4033 : _T_216;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_17_inst <= _T_44010 & _T_25 ? 32'h4033 : _T_4 ? (_T_97 | _T_242 ? 32'h4033 : _T_217) : _T_242 ?
                                32'h4033 : _T_217;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_18_inst <= _T_44010 & _T_26 ? 32'h4033 : _T_4 ? (_T_98 | _T_243 ? 32'h4033 : _T_218) : _T_243 ?
                                32'h4033 : _T_218;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_19_inst <= _T_44010 & _T_27 ? 32'h4033 : _T_4 ? (_T_99 | _T_244 ? 32'h4033 : _T_219) : _T_244 ?
                                32'h4033 : _T_219;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_20_inst <= _T_44010 & _T_28 ? 32'h4033 : _T_4 ? (_T_100 | _T_245 ? 32'h4033 : _T_220) : _T_245 ?
                                32'h4033 : _T_220;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_21_inst <= _T_44010 & _T_29 ? 32'h4033 : _T_4 ? (_T_101 | _T_246 ? 32'h4033 : _T_221) : _T_246 ?
                                32'h4033 : _T_221;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_22_inst <= _T_44010 & _T_30 ? 32'h4033 : _T_4 ? (_T_102 | _T_247 ? 32'h4033 : _T_222) : _T_247 ?
                                32'h4033 : _T_222;	// rob.scala:357:33, :487:35, :515:33, :519:33
    T_38110_23_inst <= _T_44010 & _T_31 ? 32'h4033 : _T_4 ? (_T_103 | _T_248 ? 32'h4033 : _T_223) : _T_248 ?
                                32'h4033 : _T_223;	// rob.scala:357:33, :487:35, :515:33, :519:33
    `ifndef SYNTHESIS	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_44285)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_44285)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_44297)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_44297)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
      if (`PRINTF_COND_ & ~_T_44489)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_44489)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_44501)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_44501)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
    `endif
    T_38110_0_debug_wdata <= _T_44507 & _T_176 ? io_debug_wb_wdata_2 : _T_44303 & _T_152 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_128 ? io_debug_wb_wdata_0 : ~io_dis_valids_1 | |rob_tail ?
                                T_38110_0_debug_wdata : io_dis_uops_1_debug_wdata;	// rob.scala:192:32, :347:34, :350:34, :531:53
    T_38110_1_debug_wdata <= _T_44507 & _T_177 ? io_debug_wb_wdata_2 : _T_44303 & _T_153 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_129 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_9 ?
                                io_dis_uops_1_debug_wdata : T_38110_1_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_2_debug_wdata <= _T_44507 & _T_178 ? io_debug_wb_wdata_2 : _T_44303 & _T_154 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_130 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_10 ?
                                io_dis_uops_1_debug_wdata : T_38110_2_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_3_debug_wdata <= _T_44507 & _T_179 ? io_debug_wb_wdata_2 : _T_44303 & _T_155 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_131 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_11 ?
                                io_dis_uops_1_debug_wdata : T_38110_3_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_4_debug_wdata <= _T_44507 & _T_180 ? io_debug_wb_wdata_2 : _T_44303 & _T_156 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_132 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_12 ?
                                io_dis_uops_1_debug_wdata : T_38110_4_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_5_debug_wdata <= _T_44507 & _T_181 ? io_debug_wb_wdata_2 : _T_44303 & _T_157 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_133 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_13 ?
                                io_dis_uops_1_debug_wdata : T_38110_5_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_6_debug_wdata <= _T_44507 & _T_182 ? io_debug_wb_wdata_2 : _T_44303 & _T_158 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_134 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_14 ?
                                io_dis_uops_1_debug_wdata : T_38110_6_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_7_debug_wdata <= _T_44507 & _T_183 ? io_debug_wb_wdata_2 : _T_44303 & _T_159 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_135 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_15 ?
                                io_dis_uops_1_debug_wdata : T_38110_7_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_8_debug_wdata <= _T_44507 & _T_184 ? io_debug_wb_wdata_2 : _T_44303 & _T_160 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_136 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_16 ?
                                io_dis_uops_1_debug_wdata : T_38110_8_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_9_debug_wdata <= _T_44507 & _T_185 ? io_debug_wb_wdata_2 : _T_44303 & _T_161 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_137 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_17 ?
                                io_dis_uops_1_debug_wdata : T_38110_9_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_10_debug_wdata <= _T_44507 & _T_186 ? io_debug_wb_wdata_2 : _T_44303 & _T_162 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_138 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_18 ?
                                io_dis_uops_1_debug_wdata : T_38110_10_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_11_debug_wdata <= _T_44507 & _T_187 ? io_debug_wb_wdata_2 : _T_44303 & _T_163 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_139 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_19 ?
                                io_dis_uops_1_debug_wdata : T_38110_11_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_12_debug_wdata <= _T_44507 & _T_188 ? io_debug_wb_wdata_2 : _T_44303 & _T_164 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_140 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_20 ?
                                io_dis_uops_1_debug_wdata : T_38110_12_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_13_debug_wdata <= _T_44507 & _T_189 ? io_debug_wb_wdata_2 : _T_44303 & _T_165 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_141 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_21 ?
                                io_dis_uops_1_debug_wdata : T_38110_13_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_14_debug_wdata <= _T_44507 & _T_190 ? io_debug_wb_wdata_2 : _T_44303 & _T_166 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_142 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_22 ?
                                io_dis_uops_1_debug_wdata : T_38110_14_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_15_debug_wdata <= _T_44507 & _T_191 ? io_debug_wb_wdata_2 : _T_44303 & _T_167 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_143 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_23 ?
                                io_dis_uops_1_debug_wdata : T_38110_15_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_16_debug_wdata <= _T_44507 & _T_192 ? io_debug_wb_wdata_2 : _T_44303 & _T_168 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_144 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_24 ?
                                io_dis_uops_1_debug_wdata : T_38110_16_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_17_debug_wdata <= _T_44507 & _T_193 ? io_debug_wb_wdata_2 : _T_44303 & _T_169 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_145 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_25 ?
                                io_dis_uops_1_debug_wdata : T_38110_17_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_18_debug_wdata <= _T_44507 & _T_194 ? io_debug_wb_wdata_2 : _T_44303 & _T_170 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_146 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_26 ?
                                io_dis_uops_1_debug_wdata : T_38110_18_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_19_debug_wdata <= _T_44507 & _T_195 ? io_debug_wb_wdata_2 : _T_44303 & _T_171 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_147 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_27 ?
                                io_dis_uops_1_debug_wdata : T_38110_19_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_20_debug_wdata <= _T_44507 & _T_196 ? io_debug_wb_wdata_2 : _T_44303 & _T_172 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_148 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_28 ?
                                io_dis_uops_1_debug_wdata : T_38110_20_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_21_debug_wdata <= _T_44507 & _T_197 ? io_debug_wb_wdata_2 : _T_44303 & _T_173 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_149 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_29 ?
                                io_dis_uops_1_debug_wdata : T_38110_21_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_22_debug_wdata <= _T_44507 & _T_198 ? io_debug_wb_wdata_2 : _T_44303 & _T_174 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_150 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_30 ?
                                io_dis_uops_1_debug_wdata : T_38110_22_debug_wdata;	// rob.scala:350:34, :531:53
    T_38110_23_debug_wdata <= _T_44507 & _T_199 ? io_debug_wb_wdata_2 : _T_44303 & _T_175 ? io_debug_wb_wdata_1 :
                                _T_44099 & _T_151 ? io_debug_wb_wdata_0 : io_dis_valids_1 & _T_31 ?
                                io_dis_uops_1_debug_wdata : T_38110_23_debug_wdata;	// rob.scala:350:34, :531:53
    `ifndef SYNTHESIS	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_44693)	// rob.scala:535:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to an invalid ROB entry.\n    at rob.scala:535 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:535:17
      if (`STOP_COND_ & ~_T_44693)	// rob.scala:535:17
        $fatal;	// rob.scala:535:17
      if (`PRINTF_COND_ & ~_T_44705)	// rob.scala:535:17, :538:17
        $fwrite(32'h80000002, "Assertion failed: [ROB] writeback occurred to the wrong pdst.\n    at rob.scala:538 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:538:17
      if (`STOP_COND_ & ~_T_44705)	// rob.scala:535:17, :538:17
        $fatal;	// rob.scala:538:17
    `endif
    T_47576 <= _T_47568 & _T_47569;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2941:13, rob.scala:601:48
    T_47616 <= _T_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:2979:13
    `ifndef SYNTHESIS	// rob.scala:630:14
      if (`PRINTF_COND_ & ~_T_47646)	// rob.scala:630:14
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:630 assert (!(io.com_valids(w) &&\n");	// rob.scala:630:14
      if (`STOP_COND_ & ~_T_47646)	// rob.scala:630:14
        $fatal;	// rob.scala:630:14
      if (`PRINTF_COND_ & ~_T_47657)	// rob.scala:630:14, :634:14
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:634 assert (!(io.com_valids(w) &&\n");	// rob.scala:634:14
      if (`STOP_COND_ & ~_T_47657)	// rob.scala:630:14, :634:14
        $fatal;	// rob.scala:634:14
      if (`PRINTF_COND_ & ~_T_47675)	// rob.scala:630:14
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:630 assert (!(io.com_valids(w) &&\n");	// rob.scala:630:14
      if (`STOP_COND_ & ~_T_47675)	// rob.scala:630:14
        $fatal;	// rob.scala:630:14
      if (`PRINTF_COND_ & ~_T_47686)	// rob.scala:630:14, :634:14
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:634 assert (!(io.com_valids(w) &&\n");	// rob.scala:634:14
      if (`STOP_COND_ & ~_T_47686)	// rob.scala:630:14, :634:14
        $fatal;	// rob.scala:634:14
    `endif
    if (_T_47875) begin	// rob.scala:681:26
      r_xcpt_badvaddr <= _T_249 ? io_dis_uops_0_pc + {37'h0, ~_T_47869, 2'h0} : _T_47876 & _T_47981 ?
                                                (io_lxcpt_valid ? io_lxcpt_bits_badvaddr : io_bxcpt_bits_badvaddr) : r_xcpt_badvaddr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:12:59, rob.scala:672:{37,43}, :677:40, :682:{26,47}, util.scala:114:43
      r_xcpt_uop_valid <= _T_249 ? (_T_47869 ? io_dis_uops_0_valid : io_dis_uops_1_valid) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_valid : io_bxcpt_bits_uop_valid) : r_xcpt_uop_valid;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_iw_state <= _T_249 ? (_T_47869 ? io_dis_uops_0_iw_state : io_dis_uops_1_iw_state) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_iw_state : io_bxcpt_bits_uop_iw_state) :
                                                r_xcpt_uop_iw_state;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_uopc <= _T_249 ? (_T_47869 ? io_dis_uops_0_uopc : io_dis_uops_1_uopc) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_uopc : io_bxcpt_bits_uop_uopc) : r_xcpt_uop_uopc;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_inst <= _T_249 ? (_T_47869 ? io_dis_uops_0_inst : io_dis_uops_1_inst) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_inst : io_bxcpt_bits_uop_inst) : r_xcpt_uop_inst;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_pc <= _T_249 ? (_T_47869 ? io_dis_uops_0_pc : io_dis_uops_1_pc) : _T_47876 & _T_47981 ? (_T_47887
                                                ? io_lxcpt_bits_uop_pc : io_bxcpt_bits_uop_pc) : r_xcpt_uop_pc;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_fu_code <= _T_249 ? (_T_47869 ? io_dis_uops_0_fu_code : io_dis_uops_1_fu_code) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_fu_code : io_bxcpt_bits_uop_fu_code) : r_xcpt_uop_fu_code;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_br_type <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_br_type : io_dis_uops_1_ctrl_br_type) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_br_type : io_bxcpt_bits_uop_ctrl_br_type) :
                                                r_xcpt_uop_ctrl_br_type;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_op1_sel <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_op1_sel : io_dis_uops_1_ctrl_op1_sel) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_op1_sel : io_bxcpt_bits_uop_ctrl_op1_sel) :
                                                r_xcpt_uop_ctrl_op1_sel;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_op2_sel <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_op2_sel : io_dis_uops_1_ctrl_op2_sel) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_op2_sel : io_bxcpt_bits_uop_ctrl_op2_sel) :
                                                r_xcpt_uop_ctrl_op2_sel;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_imm_sel <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_imm_sel : io_dis_uops_1_ctrl_imm_sel) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_imm_sel : io_bxcpt_bits_uop_ctrl_imm_sel) :
                                                r_xcpt_uop_ctrl_imm_sel;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_op_fcn <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_op_fcn : io_dis_uops_1_ctrl_op_fcn) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_op_fcn : io_bxcpt_bits_uop_ctrl_op_fcn) :
                                                r_xcpt_uop_ctrl_op_fcn;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_fcn_dw <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_fcn_dw : io_dis_uops_1_ctrl_fcn_dw) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_fcn_dw : io_bxcpt_bits_uop_ctrl_fcn_dw) :
                                                r_xcpt_uop_ctrl_fcn_dw;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_rf_wen <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_rf_wen : io_dis_uops_1_ctrl_rf_wen) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_rf_wen : io_bxcpt_bits_uop_ctrl_rf_wen) :
                                                r_xcpt_uop_ctrl_rf_wen;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_csr_cmd <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_csr_cmd : io_dis_uops_1_ctrl_csr_cmd) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_csr_cmd : io_bxcpt_bits_uop_ctrl_csr_cmd) :
                                                r_xcpt_uop_ctrl_csr_cmd;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_is_load <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_is_load : io_dis_uops_1_ctrl_is_load) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_is_load : io_bxcpt_bits_uop_ctrl_is_load) :
                                                r_xcpt_uop_ctrl_is_load;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_is_sta <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_is_sta : io_dis_uops_1_ctrl_is_sta) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_is_sta : io_bxcpt_bits_uop_ctrl_is_sta) :
                                                r_xcpt_uop_ctrl_is_sta;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ctrl_is_std <= _T_249 ? (_T_47869 ? io_dis_uops_0_ctrl_is_std : io_dis_uops_1_ctrl_is_std) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_ctrl_is_std : io_bxcpt_bits_uop_ctrl_is_std) :
                                                r_xcpt_uop_ctrl_is_std;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_wakeup_delay <= _T_249 ? (_T_47869 ? io_dis_uops_0_wakeup_delay : io_dis_uops_1_wakeup_delay) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_wakeup_delay : io_bxcpt_bits_uop_wakeup_delay) :
                                                r_xcpt_uop_wakeup_delay;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_allocate_brtag <= _T_249 ? (_T_47869 ? io_dis_uops_0_allocate_brtag : io_dis_uops_1_allocate_brtag) :
                                                _T_47876 & _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_allocate_brtag :
                                                io_bxcpt_bits_uop_allocate_brtag) : r_xcpt_uop_allocate_brtag;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_br_or_jmp <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_br_or_jmp : io_dis_uops_1_is_br_or_jmp) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_is_br_or_jmp : io_bxcpt_bits_uop_is_br_or_jmp) :
                                                r_xcpt_uop_is_br_or_jmp;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_jump <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_jump : io_dis_uops_1_is_jump) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_jump : io_bxcpt_bits_uop_is_jump) : r_xcpt_uop_is_jump;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_jal <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_jal : io_dis_uops_1_is_jal) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_jal : io_bxcpt_bits_uop_is_jal) : r_xcpt_uop_is_jal;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_ret <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_ret : io_dis_uops_1_is_ret) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_ret : io_bxcpt_bits_uop_is_ret) : r_xcpt_uop_is_ret;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_call <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_call : io_dis_uops_1_is_call) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_call : io_bxcpt_bits_uop_is_call) : r_xcpt_uop_is_call;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_tag <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_tag : io_dis_uops_1_br_tag) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_br_tag : io_bxcpt_bits_uop_br_tag) : r_xcpt_uop_br_tag;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_prediction_bpd_predict_val <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_prediction_bpd_predict_val :
                                                io_dis_uops_1_br_prediction_bpd_predict_val) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_br_prediction_bpd_predict_val :
                                                io_bxcpt_bits_uop_br_prediction_bpd_predict_val) : r_xcpt_uop_br_prediction_bpd_predict_val;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_prediction_bpd_predict_taken <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_prediction_bpd_predict_taken :
                                                io_dis_uops_1_br_prediction_bpd_predict_taken) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_br_prediction_bpd_predict_taken :
                                                io_bxcpt_bits_uop_br_prediction_bpd_predict_taken) :
                                                r_xcpt_uop_br_prediction_bpd_predict_taken;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_prediction_btb_hit <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_prediction_btb_hit :
                                                io_dis_uops_1_br_prediction_btb_hit) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_br_prediction_btb_hit : io_bxcpt_bits_uop_br_prediction_btb_hit) :
                                                r_xcpt_uop_br_prediction_btb_hit;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_prediction_btb_predicted <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_prediction_btb_predicted :
                                                io_dis_uops_1_br_prediction_btb_predicted) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_br_prediction_btb_predicted :
                                                io_bxcpt_bits_uop_br_prediction_btb_predicted) : r_xcpt_uop_br_prediction_btb_predicted;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_br_prediction_is_br_or_jalr <= _T_249 ? (_T_47869 ? io_dis_uops_0_br_prediction_is_br_or_jalr :
                                                io_dis_uops_1_br_prediction_is_br_or_jalr) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_br_prediction_is_br_or_jalr :
                                                io_bxcpt_bits_uop_br_prediction_is_br_or_jalr) : r_xcpt_uop_br_prediction_is_br_or_jalr;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stat_brjmp_mispredicted <= _T_249 ? (_T_47869 ? io_dis_uops_0_stat_brjmp_mispredicted :
                                                io_dis_uops_1_stat_brjmp_mispredicted) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_stat_brjmp_mispredicted : io_bxcpt_bits_uop_stat_brjmp_mispredicted) :
                                                r_xcpt_uop_stat_brjmp_mispredicted;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stat_btb_made_pred <= _T_249 ? (_T_47869 ? io_dis_uops_0_stat_btb_made_pred : io_dis_uops_1_stat_btb_made_pred) :
                                                _T_47876 & _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_stat_btb_made_pred :
                                                io_bxcpt_bits_uop_stat_btb_made_pred) : r_xcpt_uop_stat_btb_made_pred;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stat_btb_mispredicted <= _T_249 ? (_T_47869 ? io_dis_uops_0_stat_btb_mispredicted :
                                                io_dis_uops_1_stat_btb_mispredicted) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_stat_btb_mispredicted : io_bxcpt_bits_uop_stat_btb_mispredicted) :
                                                r_xcpt_uop_stat_btb_mispredicted;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stat_bpd_made_pred <= _T_249 ? (_T_47869 ? io_dis_uops_0_stat_bpd_made_pred : io_dis_uops_1_stat_bpd_made_pred) :
                                                _T_47876 & _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_stat_bpd_made_pred :
                                                io_bxcpt_bits_uop_stat_bpd_made_pred) : r_xcpt_uop_stat_bpd_made_pred;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stat_bpd_mispredicted <= _T_249 ? (_T_47869 ? io_dis_uops_0_stat_bpd_mispredicted :
                                                io_dis_uops_1_stat_bpd_mispredicted) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_stat_bpd_mispredicted : io_bxcpt_bits_uop_stat_bpd_mispredicted) :
                                                r_xcpt_uop_stat_bpd_mispredicted;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_fetch_pc_lob <= _T_249 ? (_T_47869 ? io_dis_uops_0_fetch_pc_lob : io_dis_uops_1_fetch_pc_lob) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_fetch_pc_lob : io_bxcpt_bits_uop_fetch_pc_lob) :
                                                r_xcpt_uop_fetch_pc_lob;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_imm_packed <= _T_249 ? (_T_47869 ? io_dis_uops_0_imm_packed : io_dis_uops_1_imm_packed) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_imm_packed : io_bxcpt_bits_uop_imm_packed) :
                                                r_xcpt_uop_imm_packed;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_csr_addr <= _T_249 ? (_T_47869 ? io_dis_uops_0_csr_addr : io_dis_uops_1_csr_addr) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_csr_addr : io_bxcpt_bits_uop_csr_addr) :
                                                r_xcpt_uop_csr_addr;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_rob_idx <= _T_249 ? (_T_47869 ? io_dis_uops_0_rob_idx : io_dis_uops_1_rob_idx) : _T_47876 & _T_47981 ?
                                                _T_47888_rob_idx : r_xcpt_uop_rob_idx;	// rob.scala:650:80, :670:37, :681:26, :686:23
      r_xcpt_uop_ldq_idx <= _T_249 ? (_T_47869 ? io_dis_uops_0_ldq_idx : io_dis_uops_1_ldq_idx) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_ldq_idx : io_bxcpt_bits_uop_ldq_idx) : r_xcpt_uop_ldq_idx;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stq_idx <= _T_249 ? (_T_47869 ? io_dis_uops_0_stq_idx : io_dis_uops_1_stq_idx) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_stq_idx : io_bxcpt_bits_uop_stq_idx) : r_xcpt_uop_stq_idx;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_brob_idx <= _T_249 ? (_T_47869 ? io_dis_uops_0_brob_idx : io_dis_uops_1_brob_idx) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_brob_idx : io_bxcpt_bits_uop_brob_idx) :
                                                r_xcpt_uop_brob_idx;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_pdst <= _T_249 ? (_T_47869 ? io_dis_uops_0_pdst : io_dis_uops_1_pdst) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_pdst : io_bxcpt_bits_uop_pdst) : r_xcpt_uop_pdst;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_pop1 <= _T_249 ? (_T_47869 ? io_dis_uops_0_pop1 : io_dis_uops_1_pop1) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_pop1 : io_bxcpt_bits_uop_pop1) : r_xcpt_uop_pop1;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_pop2 <= _T_249 ? (_T_47869 ? io_dis_uops_0_pop2 : io_dis_uops_1_pop2) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_pop2 : io_bxcpt_bits_uop_pop2) : r_xcpt_uop_pop2;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_pop3 <= _T_249 ? (_T_47869 ? io_dis_uops_0_pop3 : io_dis_uops_1_pop3) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_pop3 : io_bxcpt_bits_uop_pop3) : r_xcpt_uop_pop3;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_prs1_busy <= _T_249 ? (_T_47869 ? io_dis_uops_0_prs1_busy : io_dis_uops_1_prs1_busy) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_prs1_busy : io_bxcpt_bits_uop_prs1_busy) :
                                                r_xcpt_uop_prs1_busy;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_prs2_busy <= _T_249 ? (_T_47869 ? io_dis_uops_0_prs2_busy : io_dis_uops_1_prs2_busy) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_prs2_busy : io_bxcpt_bits_uop_prs2_busy) :
                                                r_xcpt_uop_prs2_busy;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_prs3_busy <= _T_249 ? (_T_47869 ? io_dis_uops_0_prs3_busy : io_dis_uops_1_prs3_busy) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_prs3_busy : io_bxcpt_bits_uop_prs3_busy) :
                                                r_xcpt_uop_prs3_busy;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_stale_pdst <= _T_249 ? (_T_47869 ? io_dis_uops_0_stale_pdst : io_dis_uops_1_stale_pdst) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_stale_pdst : io_bxcpt_bits_uop_stale_pdst) :
                                                r_xcpt_uop_stale_pdst;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_exception <= _T_249 ? (_T_47869 ? io_dis_uops_0_exception : io_dis_uops_1_exception) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_exception : io_bxcpt_bits_uop_exception) :
                                                r_xcpt_uop_exception;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_exc_cause <= _T_249 ? (_T_47869 ? io_dis_uops_0_exc_cause : io_dis_uops_1_exc_cause) : _T_47876 &
                                                _T_47981 ? {60'h0, io_lxcpt_valid ? io_lxcpt_bits_cause : io_bxcpt_bits_cause} :
                                                r_xcpt_uop_exc_cause;	// rob.scala:594:45, :597:24, :671:{37,43}, :681:26, :686:23
      r_xcpt_uop_bypassable <= _T_249 ? (_T_47869 ? io_dis_uops_0_bypassable : io_dis_uops_1_bypassable) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_bypassable : io_bxcpt_bits_uop_bypassable) :
                                                r_xcpt_uop_bypassable;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_mem_cmd <= _T_249 ? (_T_47869 ? io_dis_uops_0_mem_cmd : io_dis_uops_1_mem_cmd) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_mem_cmd : io_bxcpt_bits_uop_mem_cmd) : r_xcpt_uop_mem_cmd;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_mem_typ <= _T_249 ? (_T_47869 ? io_dis_uops_0_mem_typ : io_dis_uops_1_mem_typ) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_mem_typ : io_bxcpt_bits_uop_mem_typ) : r_xcpt_uop_mem_typ;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_fence <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_fence : io_dis_uops_1_is_fence) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_is_fence : io_bxcpt_bits_uop_is_fence) :
                                                r_xcpt_uop_is_fence;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_fencei <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_fencei : io_dis_uops_1_is_fencei) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_is_fencei : io_bxcpt_bits_uop_is_fencei) :
                                                r_xcpt_uop_is_fencei;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_store <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_store : io_dis_uops_1_is_store) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_is_store : io_bxcpt_bits_uop_is_store) :
                                                r_xcpt_uop_is_store;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_amo <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_amo : io_dis_uops_1_is_amo) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_amo : io_bxcpt_bits_uop_is_amo) : r_xcpt_uop_is_amo;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_load <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_load : io_dis_uops_1_is_load) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_is_load : io_bxcpt_bits_uop_is_load) : r_xcpt_uop_is_load;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_is_unique <= _T_249 ? (_T_47869 ? io_dis_uops_0_is_unique : io_dis_uops_1_is_unique) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_is_unique : io_bxcpt_bits_uop_is_unique) :
                                                r_xcpt_uop_is_unique;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_flush_on_commit <= _T_249 ? (_T_47869 ? io_dis_uops_0_flush_on_commit : io_dis_uops_1_flush_on_commit) :
                                                _T_47876 & _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_flush_on_commit :
                                                io_bxcpt_bits_uop_flush_on_commit) : r_xcpt_uop_flush_on_commit;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ldst <= _T_249 ? (_T_47869 ? io_dis_uops_0_ldst : io_dis_uops_1_ldst) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_ldst : io_bxcpt_bits_uop_ldst) : r_xcpt_uop_ldst;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_lrs1 <= _T_249 ? (_T_47869 ? io_dis_uops_0_lrs1 : io_dis_uops_1_lrs1) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_lrs1 : io_bxcpt_bits_uop_lrs1) : r_xcpt_uop_lrs1;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_lrs2 <= _T_249 ? (_T_47869 ? io_dis_uops_0_lrs2 : io_dis_uops_1_lrs2) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_lrs2 : io_bxcpt_bits_uop_lrs2) : r_xcpt_uop_lrs2;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_lrs3 <= _T_249 ? (_T_47869 ? io_dis_uops_0_lrs3 : io_dis_uops_1_lrs3) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_lrs3 : io_bxcpt_bits_uop_lrs3) : r_xcpt_uop_lrs3;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_ldst_val <= _T_249 ? (_T_47869 ? io_dis_uops_0_ldst_val : io_dis_uops_1_ldst_val) : _T_47876 & _T_47981
                                                ? (_T_47887 ? io_lxcpt_bits_uop_ldst_val : io_bxcpt_bits_uop_ldst_val) :
                                                r_xcpt_uop_ldst_val;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_dst_rtype <= _T_249 ? (_T_47869 ? io_dis_uops_0_dst_rtype : io_dis_uops_1_dst_rtype) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_dst_rtype : io_bxcpt_bits_uop_dst_rtype) :
                                                r_xcpt_uop_dst_rtype;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_lrs1_rtype <= _T_249 ? (_T_47869 ? io_dis_uops_0_lrs1_rtype : io_dis_uops_1_lrs1_rtype) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_lrs1_rtype : io_bxcpt_bits_uop_lrs1_rtype) :
                                                r_xcpt_uop_lrs1_rtype;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_lrs2_rtype <= _T_249 ? (_T_47869 ? io_dis_uops_0_lrs2_rtype : io_dis_uops_1_lrs2_rtype) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_lrs2_rtype : io_bxcpt_bits_uop_lrs2_rtype) :
                                                r_xcpt_uop_lrs2_rtype;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_frs3_en <= _T_249 ? (_T_47869 ? io_dis_uops_0_frs3_en : io_dis_uops_1_frs3_en) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_frs3_en : io_bxcpt_bits_uop_frs3_en) : r_xcpt_uop_frs3_en;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_fp_val <= _T_249 ? (_T_47869 ? io_dis_uops_0_fp_val : io_dis_uops_1_fp_val) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_fp_val : io_bxcpt_bits_uop_fp_val) : r_xcpt_uop_fp_val;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_fp_single <= _T_249 ? (_T_47869 ? io_dis_uops_0_fp_single : io_dis_uops_1_fp_single) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_fp_single : io_bxcpt_bits_uop_fp_single) :
                                                r_xcpt_uop_fp_single;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_xcpt_if <= _T_249 ? (_T_47869 ? io_dis_uops_0_xcpt_if : io_dis_uops_1_xcpt_if) : _T_47876 & _T_47981 ?
                                                (_T_47887 ? io_lxcpt_bits_uop_xcpt_if : io_bxcpt_bits_uop_xcpt_if) : r_xcpt_uop_xcpt_if;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_replay_if <= _T_249 ? (_T_47869 ? io_dis_uops_0_replay_if : io_dis_uops_1_replay_if) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_replay_if : io_bxcpt_bits_uop_replay_if) :
                                                r_xcpt_uop_replay_if;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_debug_wdata <= _T_249 ? (_T_47869 ? io_dis_uops_0_debug_wdata : io_dis_uops_1_debug_wdata) : _T_47876 &
                                                _T_47981 ? (_T_47887 ? io_lxcpt_bits_uop_debug_wdata : io_bxcpt_bits_uop_debug_wdata) :
                                                r_xcpt_uop_debug_wdata;	// rob.scala:666:32, :670:37, :681:26, :686:23
      r_xcpt_uop_debug_events_fetch_seq <= _T_249 ? (_T_47869 ? io_dis_uops_0_debug_events_fetch_seq :
                                                io_dis_uops_1_debug_events_fetch_seq) : _T_47876 & _T_47981 ? (_T_47887 ?
                                                io_lxcpt_bits_uop_debug_events_fetch_seq : io_bxcpt_bits_uop_debug_events_fetch_seq) :
                                                r_xcpt_uop_debug_events_fetch_seq;	// rob.scala:666:32, :670:37, :681:26, :686:23
    end
    r_xcpt_uop_br_mask <= ({8{~io_brinfo_valid}} | ~io_brinfo_mask) & _T_250;	// rob.scala:687:23, util.scala:32:{17,47}
    `ifndef SYNTHESIS	// rob.scala:693:11
      if (`PRINTF_COND_ & ~_T_48103)	// rob.scala:693:11
        $fwrite(32'h80000002, "Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:693 assert (!(exception_thrown && !io.cxcpt.valid && !r_xcpt_val),\n");	// rob.scala:693:11
      if (`STOP_COND_ & ~_T_48103)	// rob.scala:693:11
        $fatal;	// rob.scala:693:11
      if (`PRINTF_COND_ & ~_T_48109)	// rob.scala:693:11, :696:11
        $fwrite(32'h80000002, "Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:696 assert (!(io.empty && r_xcpt_val),\n");	// rob.scala:696:11
      if (`STOP_COND_ & ~_T_48109)	// rob.scala:693:11, :696:11
        $fatal;	// rob.scala:696:11
      if (`PRINTF_COND_ & ~_T_48118)	// rob.scala:693:11, :699:11
        $fwrite(32'h80000002, "Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:699 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");	// rob.scala:699:11
      if (`STOP_COND_ & ~_T_48118)	// rob.scala:693:11, :699:11
        $fatal;	// rob.scala:699:11
      if (`PRINTF_COND_ & ~reset) begin	// rob.scala:693:11, :945:13, :1061:16
        $fwrite(32'h80000002, "  RobXcpt[%c%x r:%d b:%x bva:0x%x]\n", r_xcpt_val ? 8'h45 : 8'h2D, r_xcpt_uop_exc_cause, r_xcpt_uop_rob_idx, r_xcpt_uop_br_mask, _T_6);	// rob.scala:597:24, :650:80, :667:16, :670:37, :945:13, :946:18
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h0, |rob_head | |rob_tail ? (|rob_head ? (|rob_tail ? 8'h20 : 8'h54) : 8'h48) : 8'h42);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5, rob.scala:192:32, :347:34, :500:28, :967:16, :970:18, :971:18, :972:18, util.scala:76:13
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R2_data, row_metadata_has_brorjalr_R1_data, T_23706_0 ? 8'h56 : 8'h20, T_35634_0 ? 8'h56 : 8'h20, T_23710_R1_data ? 8'h42 : 8'h20, T_35638_R1_data ? 8'h42 : 8'h20, {T_23555_R1_data[28:0], 3'h0}, {T_23555_R25_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_0_inst, T_38110_0_inst, T_28311_R1_data ? 8'h45 : 8'h2D, T_40239_R1_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_185, T_26182_0_pdst, T_26182_0_br_mask, T_26182_0_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_186, T_38110_0_pdst, T_38110_0_br_mask, T_38110_0_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h1, _T_48314 & _T_48316 ? 8'h42 : _T_48314 ? 8'h48 : _T_48316 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R3_data, row_metadata_has_brorjalr_R2_data, T_23706_1 ? 8'h56 : 8'h20, T_35634_1 ? 8'h56 : 8'h20, T_23710_R2_data ? 8'h42 : 8'h20, T_35638_R2_data ? 8'h42 : 8'h20, {T_23558_R2_data[28:0], 3'h0}, {T_23558_R26_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_1_inst, T_38110_1_inst, T_28311_R2_data ? 8'h45 : 8'h2D, T_40239_R2_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_187, T_26182_1_pdst, T_26182_1_br_mask, T_26182_1_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_188, T_38110_1_pdst, T_38110_1_br_mask, T_38110_1_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h2, _T_48400 & _T_48402 ? 8'h42 : _T_48400 ? 8'h48 : _T_48402 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R4_data, row_metadata_has_brorjalr_R3_data, T_23706_2 ? 8'h56 : 8'h20, T_35634_2 ? 8'h56 : 8'h20, T_23710_R3_data ? 8'h42 : 8'h20, T_35638_R3_data ? 8'h42 : 8'h20, {T_23555_R3_data[28:0], 3'h0}, {T_23555_R27_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_2_inst, T_38110_2_inst, T_28311_R3_data ? 8'h45 : 8'h2D, T_40239_R3_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_189, T_26182_2_pdst, T_26182_2_br_mask, T_26182_2_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_190, T_38110_2_pdst, T_38110_2_br_mask, T_38110_2_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h3, _T_48486 & _T_48488 ? 8'h42 : _T_48486 ? 8'h48 : _T_48488 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R5_data, row_metadata_has_brorjalr_R4_data, T_23706_3 ? 8'h56 : 8'h20, T_35634_3 ? 8'h56 : 8'h20, T_23710_R4_data ? 8'h42 : 8'h20, T_35638_R4_data ? 8'h42 : 8'h20, {T_23558_R4_data[28:0], 3'h0}, {T_23558_R28_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_3_inst, T_38110_3_inst, T_28311_R4_data ? 8'h45 : 8'h2D, T_40239_R4_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_191, T_26182_3_pdst, T_26182_3_br_mask, T_26182_3_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_192, T_38110_3_pdst, T_38110_3_br_mask, T_38110_3_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h4, _T_48572 & _T_48574 ? 8'h42 : _T_48572 ? 8'h48 : _T_48574 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R6_data, row_metadata_has_brorjalr_R5_data, T_23706_4 ? 8'h56 : 8'h20, T_35634_4 ? 8'h56 : 8'h20, T_23710_R5_data ? 8'h42 : 8'h20, T_35638_R5_data ? 8'h42 : 8'h20, {T_23555_R5_data[28:0], 3'h0}, {T_23555_R29_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_4_inst, T_38110_4_inst, T_28311_R5_data ? 8'h45 : 8'h2D, T_40239_R5_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_193, T_26182_4_pdst, T_26182_4_br_mask, T_26182_4_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_194, T_38110_4_pdst, T_38110_4_br_mask, T_38110_4_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h5, _T_48658 & _T_48660 ? 8'h42 : _T_48658 ? 8'h48 : _T_48660 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R7_data, row_metadata_has_brorjalr_R6_data, T_23706_5 ? 8'h56 : 8'h20, T_35634_5 ? 8'h56 : 8'h20, T_23710_R6_data ? 8'h42 : 8'h20, T_35638_R6_data ? 8'h42 : 8'h20, {T_23558_R6_data[28:0], 3'h0}, {T_23558_R30_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_5_inst, T_38110_5_inst, T_28311_R6_data ? 8'h45 : 8'h2D, T_40239_R6_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_195, T_26182_5_pdst, T_26182_5_br_mask, T_26182_5_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_196, T_38110_5_pdst, T_38110_5_br_mask, T_38110_5_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h6, _T_48744 & _T_48746 ? 8'h42 : _T_48744 ? 8'h48 : _T_48746 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R8_data, row_metadata_has_brorjalr_R7_data, T_23706_6 ? 8'h56 : 8'h20, T_35634_6 ? 8'h56 : 8'h20, T_23710_R7_data ? 8'h42 : 8'h20, T_35638_R7_data ? 8'h42 : 8'h20, {T_23555_R7_data[28:0], 3'h0}, {T_23555_R31_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_6_inst, T_38110_6_inst, T_28311_R7_data ? 8'h45 : 8'h2D, T_40239_R7_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_197, T_26182_6_pdst, T_26182_6_br_mask, T_26182_6_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_198, T_38110_6_pdst, T_38110_6_br_mask, T_38110_6_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h7, _T_48830 & _T_48832 ? 8'h42 : _T_48830 ? 8'h48 : _T_48832 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R9_data, row_metadata_has_brorjalr_R8_data, T_23706_7 ? 8'h56 : 8'h20, T_35634_7 ? 8'h56 : 8'h20, T_23710_R8_data ? 8'h42 : 8'h20, T_35638_R8_data ? 8'h42 : 8'h20, {T_23558_R8_data[28:0], 3'h0}, {T_23558_R32_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_7_inst, T_38110_7_inst, T_28311_R8_data ? 8'h45 : 8'h2D, T_40239_R8_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_199, T_26182_7_pdst, T_26182_7_br_mask, T_26182_7_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_200, T_38110_7_pdst, T_38110_7_br_mask, T_38110_7_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h8, _T_48916 & _T_48918 ? 8'h42 : _T_48916 ? 8'h48 : _T_48918 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R10_data, row_metadata_has_brorjalr_R9_data, T_23706_8 ? 8'h56 : 8'h20, T_35634_8 ? 8'h56 : 8'h20, T_23710_R9_data ? 8'h42 : 8'h20, T_35638_R9_data ? 8'h42 : 8'h20, {T_23555_R9_data[28:0], 3'h0}, {T_23555_R33_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_8_inst, T_38110_8_inst, T_28311_R9_data ? 8'h45 : 8'h2D, T_40239_R9_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_201, T_26182_8_pdst, T_26182_8_br_mask, T_26182_8_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_202, T_38110_8_pdst, T_38110_8_br_mask, T_38110_8_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h9, _T_49002 & _T_49004 ? 8'h42 : _T_49002 ? 8'h48 : _T_49004 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R11_data, row_metadata_has_brorjalr_R10_data, T_23706_9 ? 8'h56 : 8'h20, T_35634_9 ? 8'h56 : 8'h20, T_23710_R10_data ? 8'h42 : 8'h20, T_35638_R10_data ? 8'h42 : 8'h20, {T_23558_R10_data[28:0], 3'h0}, {T_23558_R34_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_9_inst, T_38110_9_inst, T_28311_R10_data ? 8'h45 : 8'h2D, T_40239_R10_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_203, T_26182_9_pdst, T_26182_9_br_mask, T_26182_9_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_204, T_38110_9_pdst, T_38110_9_br_mask, T_38110_9_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hA, _T_49088 & _T_49090 ? 8'h42 : _T_49088 ? 8'h48 : _T_49090 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R12_data, row_metadata_has_brorjalr_R11_data, T_23706_10 ? 8'h56 : 8'h20, T_35634_10 ? 8'h56 : 8'h20, T_23710_R11_data ? 8'h42 : 8'h20, T_35638_R11_data ? 8'h42 : 8'h20, {T_23555_R11_data[28:0], 3'h0}, {T_23555_R35_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_10_inst, T_38110_10_inst, T_28311_R11_data ? 8'h45 : 8'h2D, T_40239_R11_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_205, T_26182_10_pdst, T_26182_10_br_mask, T_26182_10_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_206, T_38110_10_pdst, T_38110_10_br_mask, T_38110_10_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hB, _T_49174 & _T_49176 ? 8'h42 : _T_49174 ? 8'h48 : _T_49176 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R13_data, row_metadata_has_brorjalr_R12_data, T_23706_11 ? 8'h56 : 8'h20, T_35634_11 ? 8'h56 : 8'h20, T_23710_R12_data ? 8'h42 : 8'h20, T_35638_R12_data ? 8'h42 : 8'h20, {T_23558_R12_data[28:0], 3'h0}, {T_23558_R36_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_11_inst, T_38110_11_inst, T_28311_R12_data ? 8'h45 : 8'h2D, T_40239_R12_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_207, T_26182_11_pdst, T_26182_11_br_mask, T_26182_11_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_208, T_38110_11_pdst, T_38110_11_br_mask, T_38110_11_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hC, _T_49260 & _T_49262 ? 8'h42 : _T_49260 ? 8'h48 : _T_49262 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R14_data, row_metadata_has_brorjalr_R13_data, T_23706_12 ? 8'h56 : 8'h20, T_35634_12 ? 8'h56 : 8'h20, T_23710_R13_data ? 8'h42 : 8'h20, T_35638_R13_data ? 8'h42 : 8'h20, {T_23555_R13_data[28:0], 3'h0}, {T_23555_R37_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_12_inst, T_38110_12_inst, T_28311_R13_data ? 8'h45 : 8'h2D, T_40239_R13_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_209, T_26182_12_pdst, T_26182_12_br_mask, T_26182_12_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_210, T_38110_12_pdst, T_38110_12_br_mask, T_38110_12_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hD, _T_49346 & _T_49348 ? 8'h42 : _T_49346 ? 8'h48 : _T_49348 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R15_data, row_metadata_has_brorjalr_R14_data, T_23706_13 ? 8'h56 : 8'h20, T_35634_13 ? 8'h56 : 8'h20, T_23710_R14_data ? 8'h42 : 8'h20, T_35638_R14_data ? 8'h42 : 8'h20, {T_23558_R14_data[28:0], 3'h0}, {T_23558_R38_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_13_inst, T_38110_13_inst, T_28311_R14_data ? 8'h45 : 8'h2D, T_40239_R14_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_211, T_26182_13_pdst, T_26182_13_br_mask, T_26182_13_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_212, T_38110_13_pdst, T_38110_13_br_mask, T_38110_13_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hE, _T_49432 & _T_49434 ? 8'h42 : _T_49432 ? 8'h48 : _T_49434 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R16_data, row_metadata_has_brorjalr_R15_data, T_23706_14 ? 8'h56 : 8'h20, T_35634_14 ? 8'h56 : 8'h20, T_23710_R15_data ? 8'h42 : 8'h20, T_35638_R15_data ? 8'h42 : 8'h20, {T_23555_R15_data[28:0], 3'h0}, {T_23555_R39_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_14_inst, T_38110_14_inst, T_28311_R15_data ? 8'h45 : 8'h2D, T_40239_R15_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_213, T_26182_14_pdst, T_26182_14_br_mask, T_26182_14_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_214, T_38110_14_pdst, T_38110_14_br_mask, T_38110_14_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'hF, _T_49518 & _T_49520 ? 8'h42 : _T_49518 ? 8'h48 : _T_49520 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R17_data, row_metadata_has_brorjalr_R16_data, T_23706_15 ? 8'h56 : 8'h20, T_35634_15 ? 8'h56 : 8'h20, T_23710_R16_data ? 8'h42 : 8'h20, T_35638_R16_data ? 8'h42 : 8'h20, {T_23558_R16_data[28:0], 3'h0}, {T_23558_R40_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_15_inst, T_38110_15_inst, T_28311_R16_data ? 8'h45 : 8'h2D, T_40239_R16_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_215, T_26182_15_pdst, T_26182_15_br_mask, T_26182_15_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_216, T_38110_15_pdst, T_38110_15_br_mask, T_38110_15_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h10, _T_49604 & _T_49606 ? 8'h42 : _T_49604 ? 8'h48 : _T_49606 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R18_data, row_metadata_has_brorjalr_R17_data, T_23706_16 ? 8'h56 : 8'h20, T_35634_16 ? 8'h56 : 8'h20, T_23710_R17_data ? 8'h42 : 8'h20, T_35638_R17_data ? 8'h42 : 8'h20, {T_23555_R17_data[28:0], 3'h0}, {T_23555_R41_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_16_inst, T_38110_16_inst, T_28311_R17_data ? 8'h45 : 8'h2D, T_40239_R17_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_217, T_26182_16_pdst, T_26182_16_br_mask, T_26182_16_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_218, T_38110_16_pdst, T_38110_16_br_mask, T_38110_16_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h11, _T_49690 & _T_49692 ? 8'h42 : _T_49690 ? 8'h48 : _T_49692 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R19_data, row_metadata_has_brorjalr_R18_data, T_23706_17 ? 8'h56 : 8'h20, T_35634_17 ? 8'h56 : 8'h20, T_23710_R18_data ? 8'h42 : 8'h20, T_35638_R18_data ? 8'h42 : 8'h20, {T_23558_R18_data[28:0], 3'h0}, {T_23558_R42_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_17_inst, T_38110_17_inst, T_28311_R18_data ? 8'h45 : 8'h2D, T_40239_R18_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_219, T_26182_17_pdst, T_26182_17_br_mask, T_26182_17_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_220, T_38110_17_pdst, T_38110_17_br_mask, T_38110_17_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h12, _T_49776 & _T_49778 ? 8'h42 : _T_49776 ? 8'h48 : _T_49778 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R20_data, row_metadata_has_brorjalr_R19_data, T_23706_18 ? 8'h56 : 8'h20, T_35634_18 ? 8'h56 : 8'h20, T_23710_R19_data ? 8'h42 : 8'h20, T_35638_R19_data ? 8'h42 : 8'h20, {T_23555_R19_data[28:0], 3'h0}, {T_23555_R43_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_18_inst, T_38110_18_inst, T_28311_R19_data ? 8'h45 : 8'h2D, T_40239_R19_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_221, T_26182_18_pdst, T_26182_18_br_mask, T_26182_18_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_222, T_38110_18_pdst, T_38110_18_br_mask, T_38110_18_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h13, _T_49862 & _T_49864 ? 8'h42 : _T_49862 ? 8'h48 : _T_49864 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R21_data, row_metadata_has_brorjalr_R20_data, T_23706_19 ? 8'h56 : 8'h20, T_35634_19 ? 8'h56 : 8'h20, T_23710_R20_data ? 8'h42 : 8'h20, T_35638_R20_data ? 8'h42 : 8'h20, {T_23558_R20_data[28:0], 3'h0}, {T_23558_R44_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_19_inst, T_38110_19_inst, T_28311_R20_data ? 8'h45 : 8'h2D, T_40239_R20_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_223, T_26182_19_pdst, T_26182_19_br_mask, T_26182_19_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_224, T_38110_19_pdst, T_38110_19_br_mask, T_38110_19_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h14, _T_49948 & _T_49950 ? 8'h42 : _T_49948 ? 8'h48 : _T_49950 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R22_data, row_metadata_has_brorjalr_R21_data, T_23706_20 ? 8'h56 : 8'h20, T_35634_20 ? 8'h56 : 8'h20, T_23710_R21_data ? 8'h42 : 8'h20, T_35638_R21_data ? 8'h42 : 8'h20, {T_23555_R21_data[28:0], 3'h0}, {T_23555_R45_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_20_inst, T_38110_20_inst, T_28311_R21_data ? 8'h45 : 8'h2D, T_40239_R21_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_225, T_26182_20_pdst, T_26182_20_br_mask, T_26182_20_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_226, T_38110_20_pdst, T_38110_20_br_mask, T_38110_20_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h15, _T_50034 & _T_50036 ? 8'h42 : _T_50034 ? 8'h48 : _T_50036 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R23_data, row_metadata_has_brorjalr_R22_data, T_23706_21 ? 8'h56 : 8'h20, T_35634_21 ? 8'h56 : 8'h20, T_23710_R22_data ? 8'h42 : 8'h20, T_35638_R22_data ? 8'h42 : 8'h20, {T_23558_R22_data[28:0], 3'h0}, {T_23558_R46_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_21_inst, T_38110_21_inst, T_28311_R22_data ? 8'h45 : 8'h2D, T_40239_R22_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_227, T_26182_21_pdst, T_26182_21_br_mask, T_26182_21_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_228, T_38110_21_pdst, T_38110_21_br_mask, T_38110_21_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h16, _T_50120 & _T_50122 ? 8'h42 : _T_50120 ? 8'h48 : _T_50122 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R24_data, row_metadata_has_brorjalr_R23_data, T_23706_22 ? 8'h56 : 8'h20, T_35634_22 ? 8'h56 : 8'h20, T_23710_R23_data ? 8'h42 : 8'h20, T_35638_R23_data ? 8'h42 : 8'h20, {T_23555_R23_data[28:0], 3'h0}, {T_23555_R47_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_22_inst, T_38110_22_inst, T_28311_R23_data ? 8'h45 : 8'h2D, T_40239_R23_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :893:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_229, T_26182_22_pdst, T_26182_22_br_mask, T_26182_22_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_230, T_38110_22_pdst, T_38110_22_br_mask, T_38110_22_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
        $fwrite(32'h80000002, "    rob[%d] %c (", 6'h17, _T_50206 & _T_48185 ? 8'h42 : _T_50206 ? 8'h48 : _T_48185 ? 8'h54 : 8'h20);	// rob.scala:967:16, :970:{18,40}, :971:18, :972:18
        $fwrite(32'h80000002, "%d %x (%c%c)(%c%c) 0x%x %x [%cDASM(%x)][DASM(%x) ] %c,%c ", row_metadata_brob_idx_R25_data, row_metadata_has_brorjalr_R24_data, T_23706_23 ? 8'h56 : 8'h20, T_35634_23 ? 8'h56 : 8'h20, T_23710_R24_data ? 8'h42 : 8'h20, T_35638_R24_data ? 8'h42 : 8'h20, {T_23558_R24_data[28:0], 3'h0}, {T_23558_R48_data[12:0], 3'h0} + 16'h4, 8'h20, T_26182_23_inst, T_38110_23_inst, T_28311_R24_data ? 8'h45 : 8'h2D, T_40239_R24_data ? 8'h45 : 8'h2D);	// Mux.scala:31:69, rob.scala:295:35, :296:38, :335:30, :339:30, :347:34, :350:34, :554:94, :894:22, :946:18, :970:18, :972:18, :993:19, :996:21, :997:21, :998:21, :999:21, :1000:45, :1007:21, :1008:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_231, T_26182_23_pdst, T_26182_23_br_mask, T_26182_23_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "(d:%c p%d, bm:%x sdt:%d) ", casez_tmp_232, T_38110_23_pdst, T_38110_23_br_mask, T_38110_23_stale_pdst);	// rob.scala:350:34, :1047:19, :1048:21
        $fwrite(32'h80000002, "\n");	// rob.scala:1061:16
      end
    `endif
  end // always @(posedge)
  T_23555_ext T_23555 (	// rob.scala:893:22
    .R0_addr  (_io_get_pc_rob_idx_1 ? (_io_get_pc_rob_idx_5to2 == 4'hB ? 4'h0 : _io_get_pc_rob_idx_5to2 +
                4'h1) : _io_get_pc_rob_idx_5to2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5, :964:5, rob.scala:913:29, util.scala:75:28, :76:{13,35}
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (4'h8),	// rob.scala:276:51
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (4'h8),	// rob.scala:276:51
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (4'h9),	// rob.scala:487:35
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (4'h9),	// rob.scala:487:35
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (4'hA),	// rob.scala:487:35
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (4'hA),	// rob.scala:487:35
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (4'hB),	// util.scala:75:28
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (4'hB),	// util.scala:75:28
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .R25_addr (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R25_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R25_clk  (clk),
    .R26_addr (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R26_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R26_clk  (clk),
    .R27_addr (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R27_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R27_clk  (clk),
    .R28_addr (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R28_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R28_clk  (clk),
    .R29_addr (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R29_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R29_clk  (clk),
    .R30_addr (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R30_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R30_clk  (clk),
    .R31_addr (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R31_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R31_clk  (clk),
    .R32_addr (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R32_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R32_clk  (clk),
    .R33_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R33_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R33_clk  (clk),
    .R34_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R34_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R34_clk  (clk),
    .R35_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R35_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R35_clk  (clk),
    .R36_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R36_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R36_clk  (clk),
    .R37_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R37_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R37_clk  (clk),
    .R38_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R38_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R38_clk  (clk),
    .R39_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R39_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R39_clk  (clk),
    .R40_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R40_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R40_clk  (clk),
    .R41_addr (4'h8),	// rob.scala:276:51
    .R41_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R41_clk  (clk),
    .R42_addr (4'h8),	// rob.scala:276:51
    .R42_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R42_clk  (clk),
    .R43_addr (4'h9),	// rob.scala:487:35
    .R43_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R43_clk  (clk),
    .R44_addr (4'h9),	// rob.scala:487:35
    .R44_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R44_clk  (clk),
    .R45_addr (4'hA),	// rob.scala:487:35
    .R45_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R45_clk  (clk),
    .R46_addr (4'hA),	// rob.scala:487:35
    .R46_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R46_clk  (clk),
    .R47_addr (4'hB),	// util.scala:75:28
    .R47_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R47_clk  (clk),
    .R48_addr (4'hB),	// util.scala:75:28
    .R48_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R48_clk  (clk),
    .R49_addr (_rob_head_4to1),
    .R49_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R49_clk  (clk),
    .W0_addr  (_rob_tail_4to1),
    .W0_en    (_T_23559 & ~_T_23563),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:56:9, rob.scala:933:10
    .W0_clk   (clk),
    .W0_data  (_io_dis_uops_0_pc_39to3),
    .R0_data  (T_23555_R0_data),
    .R1_data  (T_23555_R1_data),
    .R2_data  (T_23555_R2_data),
    .R3_data  (T_23555_R3_data),
    .R4_data  (T_23555_R4_data),
    .R5_data  (T_23555_R5_data),
    .R6_data  (T_23555_R6_data),
    .R7_data  (T_23555_R7_data),
    .R8_data  (T_23555_R8_data),
    .R9_data  (T_23555_R9_data),
    .R10_data (T_23555_R10_data),
    .R11_data (T_23555_R11_data),
    .R12_data (T_23555_R12_data),
    .R13_data (T_23555_R13_data),
    .R14_data (T_23555_R14_data),
    .R15_data (T_23555_R15_data),
    .R16_data (T_23555_R16_data),
    .R17_data (T_23555_R17_data),
    .R18_data (T_23555_R18_data),
    .R19_data (T_23555_R19_data),
    .R20_data (T_23555_R20_data),
    .R21_data (T_23555_R21_data),
    .R22_data (T_23555_R22_data),
    .R23_data (T_23555_R23_data),
    .R24_data (T_23555_R24_data),
    .R25_data (T_23555_R25_data),
    .R26_data (T_23555_R26_data),
    .R27_data (T_23555_R27_data),
    .R28_data (T_23555_R28_data),
    .R29_data (T_23555_R29_data),
    .R30_data (T_23555_R30_data),
    .R31_data (T_23555_R31_data),
    .R32_data (T_23555_R32_data),
    .R33_data (T_23555_R33_data),
    .R34_data (T_23555_R34_data),
    .R35_data (T_23555_R35_data),
    .R36_data (T_23555_R36_data),
    .R37_data (T_23555_R37_data),
    .R38_data (T_23555_R38_data),
    .R39_data (T_23555_R39_data),
    .R40_data (T_23555_R40_data),
    .R41_data (T_23555_R41_data),
    .R42_data (T_23555_R42_data),
    .R43_data (T_23555_R43_data),
    .R44_data (T_23555_R44_data),
    .R45_data (T_23555_R45_data),
    .R46_data (T_23555_R46_data),
    .R47_data (T_23555_R47_data),
    .R48_data (T_23555_R48_data),
    .R49_data (T_23555_R49_data)
  );
  T_23555_ext T_23558 (	// rob.scala:894:22
    .R0_addr  (_io_get_pc_rob_idx_5to2),
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R1_en    (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R3_en    (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R5_en    (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R7_en    (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R9_en    (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R11_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R13_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R15_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (4'h8),	// rob.scala:276:51
    .R17_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (4'h8),	// rob.scala:276:51
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (4'h9),	// rob.scala:487:35
    .R19_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (4'h9),	// rob.scala:487:35
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (4'hA),	// rob.scala:487:35
    .R21_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (4'hA),	// rob.scala:487:35
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (4'hB),	// util.scala:75:28
    .R23_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (4'hB),	// util.scala:75:28
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .R25_addr (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R25_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R25_clk  (clk),
    .R26_addr (4'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:912:5
    .R26_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R26_clk  (clk),
    .R27_addr (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R27_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R27_clk  (clk),
    .R28_addr (4'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:964:5
    .R28_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R28_clk  (clk),
    .R29_addr (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R29_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R29_clk  (clk),
    .R30_addr (4'h2),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1016:5
    .R30_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R30_clk  (clk),
    .R31_addr (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R31_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R31_clk  (clk),
    .R32_addr (4'h3),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1068:5
    .R32_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R32_clk  (clk),
    .R33_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R33_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R33_clk  (clk),
    .R34_addr (4'h4),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1120:5
    .R34_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R34_clk  (clk),
    .R35_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R35_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R35_clk  (clk),
    .R36_addr (4'h5),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1172:5
    .R36_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R36_clk  (clk),
    .R37_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R37_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R37_clk  (clk),
    .R38_addr (4'h6),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1224:5
    .R38_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R38_clk  (clk),
    .R39_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R39_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R39_clk  (clk),
    .R40_addr (4'h7),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:1276:5
    .R40_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R40_clk  (clk),
    .R41_addr (4'h8),	// rob.scala:276:51
    .R41_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R41_clk  (clk),
    .R42_addr (4'h8),	// rob.scala:276:51
    .R42_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R42_clk  (clk),
    .R43_addr (4'h9),	// rob.scala:487:35
    .R43_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R43_clk  (clk),
    .R44_addr (4'h9),	// rob.scala:487:35
    .R44_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R44_clk  (clk),
    .R45_addr (4'hA),	// rob.scala:487:35
    .R45_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R45_clk  (clk),
    .R46_addr (4'hA),	// rob.scala:487:35
    .R46_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R46_clk  (clk),
    .R47_addr (4'hB),	// util.scala:75:28
    .R47_en   (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R47_clk  (clk),
    .R48_addr (4'hB),	// util.scala:75:28
    .R48_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R48_clk  (clk),
    .R49_addr (_rob_head_4to1),
    .R49_en   (_T_47590),
    .R49_clk  (clk),
    .W0_addr  (_rob_tail_4to1),
    .W0_en    (_T_23559 & _T_23563),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:50:9
    .W0_clk   (clk),
    .W0_data  (_io_dis_uops_0_pc_39to3),
    .R0_data  (T_23558_R0_data),
    .R1_data  (T_23558_R1_data),
    .R2_data  (T_23558_R2_data),
    .R3_data  (T_23558_R3_data),
    .R4_data  (T_23558_R4_data),
    .R5_data  (T_23558_R5_data),
    .R6_data  (T_23558_R6_data),
    .R7_data  (T_23558_R7_data),
    .R8_data  (T_23558_R8_data),
    .R9_data  (T_23558_R9_data),
    .R10_data (T_23558_R10_data),
    .R11_data (T_23558_R11_data),
    .R12_data (T_23558_R12_data),
    .R13_data (T_23558_R13_data),
    .R14_data (T_23558_R14_data),
    .R15_data (T_23558_R15_data),
    .R16_data (T_23558_R16_data),
    .R17_data (T_23558_R17_data),
    .R18_data (T_23558_R18_data),
    .R19_data (T_23558_R19_data),
    .R20_data (T_23558_R20_data),
    .R21_data (T_23558_R21_data),
    .R22_data (T_23558_R22_data),
    .R23_data (T_23558_R23_data),
    .R24_data (T_23558_R24_data),
    .R25_data (T_23558_R25_data),
    .R26_data (T_23558_R26_data),
    .R27_data (T_23558_R27_data),
    .R28_data (T_23558_R28_data),
    .R29_data (T_23558_R29_data),
    .R30_data (T_23558_R30_data),
    .R31_data (T_23558_R31_data),
    .R32_data (T_23558_R32_data),
    .R33_data (T_23558_R33_data),
    .R34_data (T_23558_R34_data),
    .R35_data (T_23558_R35_data),
    .R36_data (T_23558_R36_data),
    .R37_data (T_23558_R37_data),
    .R38_data (T_23558_R38_data),
    .R39_data (T_23558_R39_data),
    .R40_data (T_23558_R40_data),
    .R41_data (T_23558_R41_data),
    .R42_data (T_23558_R42_data),
    .R43_data (T_23558_R43_data),
    .R44_data (T_23558_R44_data),
    .R45_data (T_23558_R45_data),
    .R46_data (T_23558_R46_data),
    .R47_data (T_23558_R47_data),
    .R48_data (T_23558_R48_data),
    .R49_data (T_23558_R49_data)
  );
  row_metadata_brob_idx_ext row_metadata_brob_idx (	// rob.scala:295:35
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (_io_get_pc_rob_idx_5to1),
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h1),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h2),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h3),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h4),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h5),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h6),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h7),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h8),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'h9),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hA),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hB),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hC),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hD),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hE),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'hF),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h10),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h11),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h12),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h13),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h14),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h15),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h16),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .R25_addr (5'h17),	// rob.scala:347:34
    .R25_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R25_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (_T_23652),
    .W0_clk   (clk),
    .W0_data  (io_dis_uops_0_brob_idx),
    .R0_data  (io_brob_deallocate_bits_brob_idx),
    .R1_data  (io_get_pc_curr_brob_idx),
    .R2_data  (row_metadata_brob_idx_R2_data),
    .R3_data  (row_metadata_brob_idx_R3_data),
    .R4_data  (row_metadata_brob_idx_R4_data),
    .R5_data  (row_metadata_brob_idx_R5_data),
    .R6_data  (row_metadata_brob_idx_R6_data),
    .R7_data  (row_metadata_brob_idx_R7_data),
    .R8_data  (row_metadata_brob_idx_R8_data),
    .R9_data  (row_metadata_brob_idx_R9_data),
    .R10_data (row_metadata_brob_idx_R10_data),
    .R11_data (row_metadata_brob_idx_R11_data),
    .R12_data (row_metadata_brob_idx_R12_data),
    .R13_data (row_metadata_brob_idx_R13_data),
    .R14_data (row_metadata_brob_idx_R14_data),
    .R15_data (row_metadata_brob_idx_R15_data),
    .R16_data (row_metadata_brob_idx_R16_data),
    .R17_data (row_metadata_brob_idx_R17_data),
    .R18_data (row_metadata_brob_idx_R18_data),
    .R19_data (row_metadata_brob_idx_R19_data),
    .R20_data (row_metadata_brob_idx_R20_data),
    .R21_data (row_metadata_brob_idx_R21_data),
    .R22_data (row_metadata_brob_idx_R22_data),
    .R23_data (row_metadata_brob_idx_R23_data),
    .R24_data (row_metadata_brob_idx_R24_data),
    .R25_data (row_metadata_brob_idx_R25_data)
  );
  row_metadata_has_brorjalr_ext row_metadata_has_brorjalr (	// rob.scala:296:38
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h1),	// rob.scala:347:34
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h2),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h3),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h4),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h5),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h6),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h7),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h8),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h9),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'hA),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hB),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hC),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hD),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hE),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hF),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'h10),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h11),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h12),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h13),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h14),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h15),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h16),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h17),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (_T_23652),
    .W0_clk   (clk),
    .W0_data  (io_dis_has_br_or_jalr_in_packet),
    .W1_addr  (rob_tail),	// rob.scala:192:32
    .W1_en    (_T_23672),
    .W1_clk   (clk),
    .W1_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_data  (row_metadata_has_brorjalr_R0_data),
    .R1_data  (row_metadata_has_brorjalr_R1_data),
    .R2_data  (row_metadata_has_brorjalr_R2_data),
    .R3_data  (row_metadata_has_brorjalr_R3_data),
    .R4_data  (row_metadata_has_brorjalr_R4_data),
    .R5_data  (row_metadata_has_brorjalr_R5_data),
    .R6_data  (row_metadata_has_brorjalr_R6_data),
    .R7_data  (row_metadata_has_brorjalr_R7_data),
    .R8_data  (row_metadata_has_brorjalr_R8_data),
    .R9_data  (row_metadata_has_brorjalr_R9_data),
    .R10_data (row_metadata_has_brorjalr_R10_data),
    .R11_data (row_metadata_has_brorjalr_R11_data),
    .R12_data (row_metadata_has_brorjalr_R12_data),
    .R13_data (row_metadata_has_brorjalr_R13_data),
    .R14_data (row_metadata_has_brorjalr_R14_data),
    .R15_data (row_metadata_has_brorjalr_R15_data),
    .R16_data (row_metadata_has_brorjalr_R16_data),
    .R17_data (row_metadata_has_brorjalr_R17_data),
    .R18_data (row_metadata_has_brorjalr_R18_data),
    .R19_data (row_metadata_has_brorjalr_R19_data),
    .R20_data (row_metadata_has_brorjalr_R20_data),
    .R21_data (row_metadata_has_brorjalr_R21_data),
    .R22_data (row_metadata_has_brorjalr_R22_data),
    .R23_data (row_metadata_has_brorjalr_R23_data),
    .R24_data (row_metadata_has_brorjalr_R24_data)
  );
  T_23710_ext T_23710 (	// rob.scala:335:30
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h1),	// rob.scala:347:34
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h2),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h3),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h4),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h5),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h6),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h7),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h8),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h9),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'hA),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hB),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hC),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hD),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hE),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hF),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'h10),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h11),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h12),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h13),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h14),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h15),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h16),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h17),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (io_dis_valids_0),
    .W0_clk   (clk),
    .W0_data  (~io_dis_uops_0_is_fence & ~io_dis_uops_0_is_fencei),	// rob.scala:348:{37,62}, :349:37
    .W1_addr  (_io_wb_resps_0_bits_uop_rob_idx_5to1),
    .W1_en    (io_wb_resps_0_valid & ~_T_28590),	// rob.scala:331:55, :368:30
    .W1_clk   (clk),
    .W1_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W2_addr  (_io_wb_resps_1_bits_uop_rob_idx_5to1),
    .W2_en    (io_wb_resps_1_valid & ~_T_28598),	// rob.scala:331:55, :368:30
    .W2_clk   (clk),
    .W2_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W3_addr  (_io_wb_resps_2_bits_uop_rob_idx_5to1),
    .W3_en    (io_wb_resps_2_valid & ~_T_28606),	// rob.scala:331:55, :368:30
    .W3_clk   (clk),
    .W3_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W4_addr  (_io_lsu_clr_bsy_rob_idx_5to1),
    .W4_en    (io_lsu_clr_bsy_valid & ~_T_28612),	// rob.scala:331:55, :388:34
    .W4_clk   (clk),
    .W4_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_data  (T_23710_R0_data),
    .R1_data  (T_23710_R1_data),
    .R2_data  (T_23710_R2_data),
    .R3_data  (T_23710_R3_data),
    .R4_data  (T_23710_R4_data),
    .R5_data  (T_23710_R5_data),
    .R6_data  (T_23710_R6_data),
    .R7_data  (T_23710_R7_data),
    .R8_data  (T_23710_R8_data),
    .R9_data  (T_23710_R9_data),
    .R10_data (T_23710_R10_data),
    .R11_data (T_23710_R11_data),
    .R12_data (T_23710_R12_data),
    .R13_data (T_23710_R13_data),
    .R14_data (T_23710_R14_data),
    .R15_data (T_23710_R15_data),
    .R16_data (T_23710_R16_data),
    .R17_data (T_23710_R17_data),
    .R18_data (T_23710_R18_data),
    .R19_data (T_23710_R19_data),
    .R20_data (T_23710_R20_data),
    .R21_data (T_23710_R21_data),
    .R22_data (T_23710_R22_data),
    .R23_data (T_23710_R23_data),
    .R24_data (T_23710_R24_data)
  );
  T_28311_ext T_28311 (	// rob.scala:339:30
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h1),	// rob.scala:347:34
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h2),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h3),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h4),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h5),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h6),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h7),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h8),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h9),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'hA),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hB),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hC),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hD),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hE),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hF),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'h10),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h11),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h12),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h13),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h14),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h15),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h16),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h17),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (io_dis_valids_0),
    .W0_clk   (clk),
    .W0_data  (io_dis_uops_0_exception),
    .W1_addr  (_io_lxcpt_bits_uop_rob_idx_5to1),
    .W1_en    (io_lxcpt_valid & ~_T_29073),	// rob.scala:331:55, :425:28
    .W1_clk   (clk),
    .W1_data  (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W2_addr  (_io_bxcpt_bits_uop_rob_idx_5to1),
    .W2_en    (io_bxcpt_valid & ~_T_29081),	// rob.scala:331:55, :429:28
    .W2_clk   (clk),
    .W2_data  (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W3_addr  (_T_2),
    .W3_en    (_T_29097),
    .W3_clk   (clk),
    .W3_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_data  (T_28311_R0_data),
    .R1_data  (T_28311_R1_data),
    .R2_data  (T_28311_R2_data),
    .R3_data  (T_28311_R3_data),
    .R4_data  (T_28311_R4_data),
    .R5_data  (T_28311_R5_data),
    .R6_data  (T_28311_R6_data),
    .R7_data  (T_28311_R7_data),
    .R8_data  (T_28311_R8_data),
    .R9_data  (T_28311_R9_data),
    .R10_data (T_28311_R10_data),
    .R11_data (T_28311_R11_data),
    .R12_data (T_28311_R12_data),
    .R13_data (T_28311_R13_data),
    .R14_data (T_28311_R14_data),
    .R15_data (T_28311_R15_data),
    .R16_data (T_28311_R16_data),
    .R17_data (T_28311_R17_data),
    .R18_data (T_28311_R18_data),
    .R19_data (T_28311_R19_data),
    .R20_data (T_28311_R20_data),
    .R21_data (T_28311_R21_data),
    .R22_data (T_28311_R22_data),
    .R23_data (T_28311_R23_data),
    .R24_data (T_28311_R24_data)
  );
  T_28314_ext T_28314 (	// rob.scala:340:30
    .R0_addr (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk  (clk),
    .W0_addr (rob_tail),	// rob.scala:192:32
    .W0_en   (io_dis_valids_0),
    .W0_clk  (clk),
    .W0_data (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .W1_addr (_io_fflags_0_bits_uop_rob_idx_5to1),
    .W1_en   (io_fflags_0_valid & ~_T_29059),	// rob.scala:331:55, :415:35
    .W1_clk  (clk),
    .W1_data (io_fflags_0_bits_flags),
    .W2_addr (_io_fflags_1_bits_uop_rob_idx_5to1),
    .W2_en   (io_fflags_1_valid & ~_T_29066),	// rob.scala:331:55, :415:35
    .W2_clk  (clk),
    .W2_data (io_fflags_1_bits_flags),
    .R0_data (T_28314_R0_data)
  );
  T_23710_ext T_35638 (	// rob.scala:335:30
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h1),	// rob.scala:347:34
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h2),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h3),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h4),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h5),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h6),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h7),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h8),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h9),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'hA),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hB),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hC),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hD),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hE),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hF),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'h10),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h11),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h12),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h13),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h14),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h15),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h16),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h17),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (io_dis_valids_1),
    .W0_clk   (clk),
    .W0_data  (~io_dis_uops_1_is_fence & ~io_dis_uops_1_is_fencei),	// rob.scala:348:{37,62}, :349:37
    .W1_addr  (_io_wb_resps_0_bits_uop_rob_idx_5to1),
    .W1_en    (io_wb_resps_0_valid & _T_28590),	// rob.scala:368:30
    .W1_clk   (clk),
    .W1_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W2_addr  (_io_wb_resps_1_bits_uop_rob_idx_5to1),
    .W2_en    (io_wb_resps_1_valid & _T_28598),	// rob.scala:368:30
    .W2_clk   (clk),
    .W2_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W3_addr  (_io_wb_resps_2_bits_uop_rob_idx_5to1),
    .W3_en    (io_wb_resps_2_valid & _T_28606),	// rob.scala:368:30
    .W3_clk   (clk),
    .W3_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W4_addr  (_io_lsu_clr_bsy_rob_idx_5to1),
    .W4_en    (io_lsu_clr_bsy_valid & _T_28612),	// rob.scala:388:34
    .W4_clk   (clk),
    .W4_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_data  (T_35638_R0_data),
    .R1_data  (T_35638_R1_data),
    .R2_data  (T_35638_R2_data),
    .R3_data  (T_35638_R3_data),
    .R4_data  (T_35638_R4_data),
    .R5_data  (T_35638_R5_data),
    .R6_data  (T_35638_R6_data),
    .R7_data  (T_35638_R7_data),
    .R8_data  (T_35638_R8_data),
    .R9_data  (T_35638_R9_data),
    .R10_data (T_35638_R10_data),
    .R11_data (T_35638_R11_data),
    .R12_data (T_35638_R12_data),
    .R13_data (T_35638_R13_data),
    .R14_data (T_35638_R14_data),
    .R15_data (T_35638_R15_data),
    .R16_data (T_35638_R16_data),
    .R17_data (T_35638_R17_data),
    .R18_data (T_35638_R18_data),
    .R19_data (T_35638_R19_data),
    .R20_data (T_35638_R20_data),
    .R21_data (T_35638_R21_data),
    .R22_data (T_35638_R22_data),
    .R23_data (T_35638_R23_data),
    .R24_data (T_35638_R24_data)
  );
  T_28311_ext T_40239 (	// rob.scala:339:30
    .R0_addr  (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk   (clk),
    .R1_addr  (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .R1_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R1_clk   (clk),
    .R2_addr  (5'h1),	// rob.scala:347:34
    .R2_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R2_clk   (clk),
    .R3_addr  (5'h2),	// rob.scala:347:34
    .R3_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R3_clk   (clk),
    .R4_addr  (5'h3),	// rob.scala:347:34
    .R4_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R4_clk   (clk),
    .R5_addr  (5'h4),	// rob.scala:347:34
    .R5_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R5_clk   (clk),
    .R6_addr  (5'h5),	// rob.scala:347:34
    .R6_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R6_clk   (clk),
    .R7_addr  (5'h6),	// rob.scala:347:34
    .R7_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R7_clk   (clk),
    .R8_addr  (5'h7),	// rob.scala:347:34
    .R8_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R8_clk   (clk),
    .R9_addr  (5'h8),	// rob.scala:347:34
    .R9_en    (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R9_clk   (clk),
    .R10_addr (5'h9),	// rob.scala:347:34
    .R10_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R10_clk  (clk),
    .R11_addr (5'hA),	// rob.scala:347:34
    .R11_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R11_clk  (clk),
    .R12_addr (5'hB),	// rob.scala:347:34
    .R12_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R12_clk  (clk),
    .R13_addr (5'hC),	// rob.scala:347:34
    .R13_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R13_clk  (clk),
    .R14_addr (5'hD),	// rob.scala:347:34
    .R14_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R14_clk  (clk),
    .R15_addr (5'hE),	// rob.scala:347:34
    .R15_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R15_clk  (clk),
    .R16_addr (5'hF),	// rob.scala:347:34
    .R16_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R16_clk  (clk),
    .R17_addr (5'h10),	// rob.scala:347:34
    .R17_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R17_clk  (clk),
    .R18_addr (5'h11),	// rob.scala:347:34
    .R18_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R18_clk  (clk),
    .R19_addr (5'h12),	// rob.scala:347:34
    .R19_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R19_clk  (clk),
    .R20_addr (5'h13),	// rob.scala:347:34
    .R20_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R20_clk  (clk),
    .R21_addr (5'h14),	// rob.scala:347:34
    .R21_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R21_clk  (clk),
    .R22_addr (5'h15),	// rob.scala:347:34
    .R22_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R22_clk  (clk),
    .R23_addr (5'h16),	// rob.scala:347:34
    .R23_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R23_clk  (clk),
    .R24_addr (5'h17),	// rob.scala:347:34
    .R24_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R24_clk  (clk),
    .W0_addr  (rob_tail),	// rob.scala:192:32
    .W0_en    (io_dis_valids_1),
    .W0_clk   (clk),
    .W0_data  (io_dis_uops_1_exception),
    .W1_addr  (_io_lxcpt_bits_uop_rob_idx_5to1),
    .W1_en    (io_lxcpt_valid & _T_29073),	// rob.scala:425:28
    .W1_clk   (clk),
    .W1_data  (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W2_addr  (_io_bxcpt_bits_uop_rob_idx_5to1),
    .W2_en    (io_bxcpt_valid & _T_29081),	// rob.scala:429:28
    .W2_clk   (clk),
    .W2_data  (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .W3_addr  (_T_2),
    .W3_en    (_T_29097),
    .W3_clk   (clk),
    .W3_data  (1'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_data  (T_40239_R0_data),
    .R1_data  (T_40239_R1_data),
    .R2_data  (T_40239_R2_data),
    .R3_data  (T_40239_R3_data),
    .R4_data  (T_40239_R4_data),
    .R5_data  (T_40239_R5_data),
    .R6_data  (T_40239_R6_data),
    .R7_data  (T_40239_R7_data),
    .R8_data  (T_40239_R8_data),
    .R9_data  (T_40239_R9_data),
    .R10_data (T_40239_R10_data),
    .R11_data (T_40239_R11_data),
    .R12_data (T_40239_R12_data),
    .R13_data (T_40239_R13_data),
    .R14_data (T_40239_R14_data),
    .R15_data (T_40239_R15_data),
    .R16_data (T_40239_R16_data),
    .R17_data (T_40239_R17_data),
    .R18_data (T_40239_R18_data),
    .R19_data (T_40239_R19_data),
    .R20_data (T_40239_R20_data),
    .R21_data (T_40239_R21_data),
    .R22_data (T_40239_R22_data),
    .R23_data (T_40239_R23_data),
    .R24_data (T_40239_R24_data)
  );
  T_28314_ext T_40242 (	// rob.scala:340:30
    .R0_addr (rob_head),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:149:5
    .R0_en   (1'h1),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
    .R0_clk  (clk),
    .W0_addr (rob_tail),	// rob.scala:192:32
    .W0_en   (io_dis_valids_1),
    .W0_clk  (clk),
    .W0_data (5'h0),	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:13:58
    .W1_addr (_io_fflags_0_bits_uop_rob_idx_5to1),
    .W1_en   (io_fflags_0_valid & _T_29059),	// rob.scala:415:35
    .W1_clk  (clk),
    .W1_data (io_fflags_0_bits_flags),
    .W2_addr (_io_fflags_1_bits_uop_rob_idx_5to1),
    .W2_en   (io_fflags_1_valid & _T_29066),	// rob.scala:415:35
    .W2_clk  (clk),
    .W2_data (io_fflags_1_bits_flags),
    .R0_data (T_40242_R0_data)
  );
  assign io_curr_rob_tail = {1'h0, rob_tail};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:192:32, util.scala:92:39
  assign io_com_valids_0 = _T_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_com_valids_1 = _T_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_com_uops_0_valid = casez_tmp_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_iw_state = casez_tmp_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_uopc = casez_tmp_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_inst = casez_tmp_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_pc = casez_tmp_8;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_fu_code = casez_tmp_9;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_br_type = casez_tmp_10;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_op1_sel = casez_tmp_11;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_op2_sel = casez_tmp_12;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_imm_sel = casez_tmp_13;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_op_fcn = casez_tmp_14;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_fcn_dw = casez_tmp_15;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_rf_wen = casez_tmp_16;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_csr_cmd = casez_tmp_17;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_is_load = casez_tmp_18;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_is_sta = casez_tmp_19;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ctrl_is_std = casez_tmp_20;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_wakeup_delay = casez_tmp_21;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_allocate_brtag = casez_tmp_22;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_br_or_jmp = casez_tmp_23;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_jump = casez_tmp_24;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_jal = casez_tmp_25;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_ret = casez_tmp_26;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_call = casez_tmp_27;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_mask = casez_tmp_28;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_tag = casez_tmp_29;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_prediction_bpd_predict_val = casez_tmp_30;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_prediction_bpd_predict_taken = casez_tmp_31;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_prediction_btb_hit = casez_tmp_32;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_prediction_btb_predicted = casez_tmp_33;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_br_prediction_is_br_or_jalr = casez_tmp_34;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stat_brjmp_mispredicted = casez_tmp_35;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stat_btb_made_pred = casez_tmp_36;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stat_btb_mispredicted = casez_tmp_37;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stat_bpd_made_pred = casez_tmp_38;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stat_bpd_mispredicted = casez_tmp_39;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_fetch_pc_lob = casez_tmp_40;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_imm_packed = casez_tmp_41;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_csr_addr = casez_tmp_42;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_rob_idx = casez_tmp_43;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ldq_idx = casez_tmp_44;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stq_idx = casez_tmp_45;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_brob_idx = casez_tmp_46;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_pdst = casez_tmp_47;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_pop1 = casez_tmp_48;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_pop2 = casez_tmp_49;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_pop3 = casez_tmp_50;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_prs1_busy = casez_tmp_51;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_prs2_busy = casez_tmp_52;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_prs3_busy = casez_tmp_53;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_stale_pdst = casez_tmp_54;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_exception = casez_tmp_55;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_exc_cause = casez_tmp_56;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_bypassable = casez_tmp_57;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_mem_cmd = casez_tmp_58;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_mem_typ = casez_tmp_59;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_fence = casez_tmp_60;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_fencei = casez_tmp_61;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_store = casez_tmp_62;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_amo = casez_tmp_63;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_load = casez_tmp_64;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_is_unique = casez_tmp_65;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_flush_on_commit = casez_tmp_66;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ldst = casez_tmp_67;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_lrs1 = casez_tmp_68;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_lrs2 = casez_tmp_69;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_lrs3 = casez_tmp_70;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_ldst_val = casez_tmp_71;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_dst_rtype = casez_tmp_72;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_lrs1_rtype = casez_tmp_73;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_lrs2_rtype = casez_tmp_74;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_frs3_en = casez_tmp_75;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_fp_val = casez_tmp_76;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_fp_single = casez_tmp_77;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_xcpt_if = casez_tmp_78;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_replay_if = casez_tmp_79;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_0_debug_wdata = casez_tmp_83;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28
  assign io_com_uops_0_debug_events_fetch_seq = casez_tmp_80;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_valid = casez_tmp_96;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_iw_state = casez_tmp_97;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_uopc = casez_tmp_98;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_inst = casez_tmp_99;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_pc = casez_tmp_100;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_fu_code = casez_tmp_101;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_br_type = casez_tmp_102;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_op1_sel = casez_tmp_103;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_op2_sel = casez_tmp_104;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_imm_sel = casez_tmp_105;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_op_fcn = casez_tmp_106;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_fcn_dw = casez_tmp_107;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_rf_wen = casez_tmp_108;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_csr_cmd = casez_tmp_109;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_is_load = casez_tmp_110;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_is_sta = casez_tmp_111;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ctrl_is_std = casez_tmp_112;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_wakeup_delay = casez_tmp_113;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_allocate_brtag = casez_tmp_114;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_br_or_jmp = casez_tmp_115;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_jump = casez_tmp_116;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_jal = casez_tmp_117;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_ret = casez_tmp_118;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_call = casez_tmp_119;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_mask = casez_tmp_120;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_tag = casez_tmp_121;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_prediction_bpd_predict_val = casez_tmp_122;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_prediction_bpd_predict_taken = casez_tmp_123;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_prediction_btb_hit = casez_tmp_124;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_prediction_btb_predicted = casez_tmp_125;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_br_prediction_is_br_or_jalr = casez_tmp_126;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stat_brjmp_mispredicted = casez_tmp_127;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stat_btb_made_pred = casez_tmp_128;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stat_btb_mispredicted = casez_tmp_129;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stat_bpd_made_pred = casez_tmp_130;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stat_bpd_mispredicted = casez_tmp_131;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_fetch_pc_lob = casez_tmp_132;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_imm_packed = casez_tmp_133;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_csr_addr = casez_tmp_134;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_rob_idx = casez_tmp_135;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ldq_idx = casez_tmp_136;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stq_idx = casez_tmp_137;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_brob_idx = casez_tmp_138;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_pdst = casez_tmp_139;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_pop1 = casez_tmp_140;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_pop2 = casez_tmp_141;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_pop3 = casez_tmp_142;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_prs1_busy = casez_tmp_143;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_prs2_busy = casez_tmp_144;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_prs3_busy = casez_tmp_145;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_stale_pdst = casez_tmp_146;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_exception = casez_tmp_147;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_exc_cause = casez_tmp_148;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_bypassable = casez_tmp_149;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_mem_cmd = casez_tmp_150;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_mem_typ = casez_tmp_151;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_fence = casez_tmp_152;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_fencei = casez_tmp_153;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_store = casez_tmp_154;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_amo = casez_tmp_155;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_load = casez_tmp_156;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_is_unique = casez_tmp_157;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_flush_on_commit = casez_tmp_158;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ldst = casez_tmp_159;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_lrs1 = casez_tmp_160;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_lrs2 = casez_tmp_161;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_lrs3 = casez_tmp_162;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_ldst_val = casez_tmp_163;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_dst_rtype = casez_tmp_164;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_lrs1_rtype = casez_tmp_165;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_lrs2_rtype = casez_tmp_166;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_frs3_en = casez_tmp_167;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_fp_val = casez_tmp_168;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_fp_single = casez_tmp_169;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_xcpt_if = casez_tmp_170;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_replay_if = casez_tmp_171;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_uops_1_debug_wdata = casez_tmp_175;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28
  assign io_com_uops_1_debug_events_fetch_seq = casez_tmp_172;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:453:59
  assign io_com_fflags_val = _T_47635 | _T_47664;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:640:44
  assign io_com_fflags = (_T_47635 ? T_28314_R0_data : 5'h0) | (_T_47664 ? T_40242_R0_data : 5'h0);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :13:58, rob.scala:340:30, :628:23, :641:40
  assign io_com_st_mask_0 = _T_3 & casez_tmp_81;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28, :869:45
  assign io_com_st_mask_1 = _T_4 & casez_tmp_173;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28, :869:45
  assign io_com_ld_mask_0 = _T_3 & casez_tmp_82;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28, :870:45
  assign io_com_ld_mask_1 = _T_4 & casez_tmp_174;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:507:28, :870:45
  assign io_com_load_is_at_rob_head = casez_tmp_2 ? casez_tmp_82 : casez_tmp_174;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:433:51, :507:28, :873:31
  assign io_com_exception = _T_47568 & ~(_T_47569 | r_xcpt_uop_exc_cause == 64'hE);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:594:77, :595:45, :596:{44,47}, :597:24
  assign io_com_exc_cause = r_xcpt_uop_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:597:24
  assign io_com_handling_exc = _T_47568;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_com_rbk_valids_0 = _T_29097 & casez_tmp_3 & (casez_tmp_72 == 2'h0 | casez_tmp_72 == 2'h1);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :12:59, rob.scala:451:58, :452:48, :453:{59,70,100}
  assign io_com_rbk_valids_1 = _T_29097 & casez_tmp_95 & (casez_tmp_164 == 2'h0 | casez_tmp_164 == 2'h1);	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :12:59, rob.scala:451:58, :452:48, :453:{59,70,100}
  assign io_com_badvaddr = {{24{r_xcpt_badvaddr[39]}}, r_xcpt_badvaddr};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, Bitwise.scala:33:12, Cat.scala:20:58, util.scala:114:43
  assign io_get_pc_curr_pc = {_io_get_pc_rob_idx_1 ? T_23558_R0_data : T_23555_R0_data, 3'h0} + {37'h0,
                io_get_pc_rob_idx[0], 2'h0};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :12:59, Mux.scala:31:69, rob.scala:227:38, :268:37, :682:47, :893:22, :894:22, :920:24
  assign io_get_pc_next_val = _rob_pc_hob_next_val | _T_23559;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:279:46
  assign io_get_pc_next_pc = _rob_pc_hob_next_val ? {_io_get_pc_rob_idx_1 ? T_23555_R0_data : T_23558_R0_data, 3'h0} +
                {37'h0, ~_T_1, 2'h0} : (io_dis_uops_0_pc & 40'hFFFFFFFFF8) + {37'h0, ~io_dis_valids_0,
                2'h0};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :12:59, Mux.scala:31:69, rob.scala:276:{51,97}, :280:28, :281:40, :509:28, :682:47, :893:22, :894:22, :921:24
  assign io_lsu_misspec = T_47576;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_flush_take_pc = _T_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_flush_pc = {_T_47590 ? T_23558_R49_data : T_23555_R49_data, 3'h0} + {37'h0, ~casez_tmp_2, 2'h0} +
                {37'h0, ~_T_47568, 2'h0};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :12:59, Mux.scala:31:69, rob.scala:433:51, :605:46, :606:86, :607:23, :682:47, :893:22, :894:22, :904:19
  assign io_flush_pipeline = T_47616;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:612:22
  assign io_flush_brob = _T_23672;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_empty = _T_48195;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
  assign io_ready = rob_state == 2'h1 & (_T_48185 ? 5'h0 : rob_tail + 5'h1) != rob_head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :13:58, :149:5, rob.scala:192:32, :347:34, :443:23, :453:100, :757:47, :764:{27,41}, util.scala:76:{13,35}
  assign io_brob_deallocate_valid = _T & row_metadata_has_brorjalr_R0_data;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:296:38, :315:56, :716:89
  assign io_debug_state = rob_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:443:23
  assign io_debug_rob_head = {1'h0, rob_head};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, :149:5, rob.scala:699:69
  assign io_debug_xcpt_val = r_xcpt_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:667:16
  assign io_debug_xcpt_uop_valid = r_xcpt_uop_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_iw_state = r_xcpt_uop_iw_state;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_uopc = r_xcpt_uop_uopc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_inst = r_xcpt_uop_inst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_pc = r_xcpt_uop_pc;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_fu_code = r_xcpt_uop_fu_code;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_br_type = r_xcpt_uop_ctrl_br_type;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_op1_sel = r_xcpt_uop_ctrl_op1_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_op2_sel = r_xcpt_uop_ctrl_op2_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_imm_sel = r_xcpt_uop_ctrl_imm_sel;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_op_fcn = r_xcpt_uop_ctrl_op_fcn;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_fcn_dw = r_xcpt_uop_ctrl_fcn_dw;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_rf_wen = r_xcpt_uop_ctrl_rf_wen;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_csr_cmd = r_xcpt_uop_ctrl_csr_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_is_load = r_xcpt_uop_ctrl_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_is_sta = r_xcpt_uop_ctrl_is_sta;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ctrl_is_std = r_xcpt_uop_ctrl_is_std;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_wakeup_delay = r_xcpt_uop_wakeup_delay;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_allocate_brtag = r_xcpt_uop_allocate_brtag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_br_or_jmp = r_xcpt_uop_is_br_or_jmp;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_jump = r_xcpt_uop_is_jump;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_jal = r_xcpt_uop_is_jal;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_ret = r_xcpt_uop_is_ret;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_call = r_xcpt_uop_is_call;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_mask = r_xcpt_uop_br_mask;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_tag = r_xcpt_uop_br_tag;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_prediction_bpd_predict_val = r_xcpt_uop_br_prediction_bpd_predict_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_prediction_bpd_predict_taken = r_xcpt_uop_br_prediction_bpd_predict_taken;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_prediction_btb_hit = r_xcpt_uop_br_prediction_btb_hit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_prediction_btb_predicted = r_xcpt_uop_br_prediction_btb_predicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_br_prediction_is_br_or_jalr = r_xcpt_uop_br_prediction_is_br_or_jalr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stat_brjmp_mispredicted = r_xcpt_uop_stat_brjmp_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stat_btb_made_pred = r_xcpt_uop_stat_btb_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stat_btb_mispredicted = r_xcpt_uop_stat_btb_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stat_bpd_made_pred = r_xcpt_uop_stat_bpd_made_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stat_bpd_mispredicted = r_xcpt_uop_stat_bpd_mispredicted;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_fetch_pc_lob = r_xcpt_uop_fetch_pc_lob;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_imm_packed = r_xcpt_uop_imm_packed;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_csr_addr = r_xcpt_uop_csr_addr;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_rob_idx = r_xcpt_uop_rob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:650:80
  assign io_debug_xcpt_uop_ldq_idx = r_xcpt_uop_ldq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stq_idx = r_xcpt_uop_stq_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_brob_idx = r_xcpt_uop_brob_idx;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_pdst = r_xcpt_uop_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_pop1 = r_xcpt_uop_pop1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_pop2 = r_xcpt_uop_pop2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_pop3 = r_xcpt_uop_pop3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_prs1_busy = r_xcpt_uop_prs1_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_prs2_busy = r_xcpt_uop_prs2_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_prs3_busy = r_xcpt_uop_prs3_busy;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_stale_pdst = r_xcpt_uop_stale_pdst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_exception = r_xcpt_uop_exception;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_exc_cause = r_xcpt_uop_exc_cause;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:597:24
  assign io_debug_xcpt_uop_bypassable = r_xcpt_uop_bypassable;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_mem_cmd = r_xcpt_uop_mem_cmd;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_mem_typ = r_xcpt_uop_mem_typ;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_fence = r_xcpt_uop_is_fence;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_fencei = r_xcpt_uop_is_fencei;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_store = r_xcpt_uop_is_store;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_amo = r_xcpt_uop_is_amo;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_load = r_xcpt_uop_is_load;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_is_unique = r_xcpt_uop_is_unique;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_flush_on_commit = r_xcpt_uop_flush_on_commit;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ldst = r_xcpt_uop_ldst;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_lrs1 = r_xcpt_uop_lrs1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_lrs2 = r_xcpt_uop_lrs2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_lrs3 = r_xcpt_uop_lrs3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_ldst_val = r_xcpt_uop_ldst_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_dst_rtype = r_xcpt_uop_dst_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_lrs1_rtype = r_xcpt_uop_lrs1_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_lrs2_rtype = r_xcpt_uop_lrs2_rtype;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_frs3_en = r_xcpt_uop_frs3_en;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_fp_val = r_xcpt_uop_fp_val;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_fp_single = r_xcpt_uop_fp_single;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_xcpt_if = r_xcpt_uop_xcpt_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_replay_if = r_xcpt_uop_replay_if;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_debug_wdata = r_xcpt_uop_debug_wdata;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_uop_debug_events_fetch_seq = r_xcpt_uop_debug_events_fetch_seq;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10, rob.scala:670:37
  assign io_debug_xcpt_badvaddr = _T_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/Rob.fir:6:10
endmodule

