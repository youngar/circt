// Standard header to adapt well known macros to our needs.
`ifdef RANDOMIZE_REG_INIT
  `define RANDOMIZE
`endif

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM {$random}
`endif

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifdef PRINTF_COND
  `define PRINTF_COND_ (`PRINTF_COND)
`else
  `define PRINTF_COND_ 1
`endif

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifdef STOP_COND
  `define STOP_COND_ (`STOP_COND)
`else
  `define STOP_COND_ 1
`endif

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifdef RANDOMIZE
  `ifdef VERILATOR
    `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
  `else
    `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
  `endif
`else
  `define INIT_RANDOM_PROLOG_
`endif

module HwachaSequencer(	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  input         clock, reset, io_op_valid,
  input  [9:0]  io_op_bits_fn_union,
  input  [63:0] io_op_bits_sreg_ss1, io_op_bits_sreg_ss2, io_op_bits_sreg_ss3,
  input  [3:0]  io_op_bits_base_vp_id,
  input         io_op_bits_base_vp_valid, io_op_bits_base_vp_scalar,
  input         io_op_bits_base_vp_pred,
  input  [7:0]  io_op_bits_base_vs1_id,
  input         io_op_bits_base_vs1_valid, io_op_bits_base_vs1_scalar,
  input         io_op_bits_base_vs1_pred,
  input  [1:0]  io_op_bits_base_vs1_prec,
  input  [7:0]  io_op_bits_base_vs2_id,
  input         io_op_bits_base_vs2_valid, io_op_bits_base_vs2_scalar,
  input         io_op_bits_base_vs2_pred,
  input  [1:0]  io_op_bits_base_vs2_prec,
  input  [7:0]  io_op_bits_base_vs3_id,
  input         io_op_bits_base_vs3_valid, io_op_bits_base_vs3_scalar,
  input         io_op_bits_base_vs3_pred,
  input  [1:0]  io_op_bits_base_vs3_prec,
  input  [7:0]  io_op_bits_base_vd_id,
  input         io_op_bits_base_vd_valid, io_op_bits_base_vd_scalar,
  input         io_op_bits_base_vd_pred,
  input  [1:0]  io_op_bits_base_vd_prec,
  input  [7:0]  io_op_bits_reg_vp_id, io_op_bits_reg_vs1_id, io_op_bits_reg_vs2_id,
  input  [7:0]  io_op_bits_reg_vs3_id, io_op_bits_reg_vd_id,
  input         io_op_bits_active_vint, io_op_bits_active_vipred,
  input         io_op_bits_active_vimul, io_op_bits_active_vidiv, io_op_bits_active_vfma,
  input         io_op_bits_active_vfdiv, io_op_bits_active_vfcmp,
  input         io_op_bits_active_vfconv, io_op_bits_active_vrpred,
  input         io_op_bits_active_vrfirst, io_op_bits_active_vamo,
  input         io_op_bits_active_vldx, io_op_bits_active_vstx, io_op_bits_active_vld,
  input         io_op_bits_active_vst, io_master_clear_0, io_master_clear_1,
  input         io_master_clear_2, io_master_clear_3, io_master_clear_4,
  input         io_master_clear_5, io_master_clear_6, io_master_clear_7, io_vf_stop,
  output        io_op_ready, io_master_state_valid_0, io_master_state_valid_1,
  output        io_master_state_valid_2, io_master_state_valid_3,
  output        io_master_state_valid_4, io_master_state_valid_5,
  output        io_master_state_valid_6, io_master_state_valid_7,
  output [9:0]  io_master_state_e_0_fn_union,
  output [63:0] io_master_state_e_0_sreg_ss1, io_master_state_e_0_sreg_ss2,
  output [63:0] io_master_state_e_0_sreg_ss3,
  output [3:0]  io_master_state_e_0_base_vp_id,
  output        io_master_state_e_0_base_vp_valid, io_master_state_e_0_base_vp_scalar,
  output        io_master_state_e_0_base_vp_pred,
  output [7:0]  io_master_state_e_0_base_vs1_id,
  output        io_master_state_e_0_base_vs1_valid, io_master_state_e_0_base_vs1_scalar,
  output        io_master_state_e_0_base_vs1_pred,
  output [1:0]  io_master_state_e_0_base_vs1_prec,
  output [7:0]  io_master_state_e_0_base_vs2_id,
  output        io_master_state_e_0_base_vs2_valid, io_master_state_e_0_base_vs2_scalar,
  output        io_master_state_e_0_base_vs2_pred,
  output [1:0]  io_master_state_e_0_base_vs2_prec,
  output [7:0]  io_master_state_e_0_base_vs3_id,
  output        io_master_state_e_0_base_vs3_valid, io_master_state_e_0_base_vs3_scalar,
  output        io_master_state_e_0_base_vs3_pred,
  output [1:0]  io_master_state_e_0_base_vs3_prec,
  output [7:0]  io_master_state_e_0_base_vd_id,
  output        io_master_state_e_0_base_vd_valid, io_master_state_e_0_base_vd_scalar,
  output        io_master_state_e_0_base_vd_pred,
  output [1:0]  io_master_state_e_0_base_vd_prec,
  output        io_master_state_e_0_rate, io_master_state_e_0_active_viu,
  output        io_master_state_e_0_active_vipu, io_master_state_e_0_active_vimu,
  output        io_master_state_e_0_active_vidu, io_master_state_e_0_active_vfmu,
  output        io_master_state_e_0_active_vfdu, io_master_state_e_0_active_vfcu,
  output        io_master_state_e_0_active_vfvu, io_master_state_e_0_active_vrpu,
  output        io_master_state_e_0_active_vrfu, io_master_state_e_0_active_vpu,
  output        io_master_state_e_0_active_vgu, io_master_state_e_0_active_vcu,
  output        io_master_state_e_0_active_vlu, io_master_state_e_0_active_vsu,
  output        io_master_state_e_0_active_vqu, io_master_state_e_0_raw_0,
  output        io_master_state_e_0_raw_1, io_master_state_e_0_raw_2,
  output        io_master_state_e_0_raw_3, io_master_state_e_0_raw_4,
  output        io_master_state_e_0_raw_5, io_master_state_e_0_raw_6,
  output        io_master_state_e_0_raw_7, io_master_state_e_0_war_0,
  output        io_master_state_e_0_war_1, io_master_state_e_0_war_2,
  output        io_master_state_e_0_war_3, io_master_state_e_0_war_4,
  output        io_master_state_e_0_war_5, io_master_state_e_0_war_6,
  output        io_master_state_e_0_war_7, io_master_state_e_0_waw_0,
  output        io_master_state_e_0_waw_1, io_master_state_e_0_waw_2,
  output        io_master_state_e_0_waw_3, io_master_state_e_0_waw_4,
  output        io_master_state_e_0_waw_5, io_master_state_e_0_waw_6,
  output        io_master_state_e_0_waw_7, io_master_state_e_0_last,
  output [1:0]  io_master_state_e_0_rports,
  output [3:0]  io_master_state_e_0_wport_sram,
  output [2:0]  io_master_state_e_0_wport_pred,
  output [9:0]  io_master_state_e_1_fn_union,
  output [63:0] io_master_state_e_1_sreg_ss1, io_master_state_e_1_sreg_ss2,
  output [63:0] io_master_state_e_1_sreg_ss3,
  output [3:0]  io_master_state_e_1_base_vp_id,
  output        io_master_state_e_1_base_vp_valid, io_master_state_e_1_base_vp_scalar,
  output        io_master_state_e_1_base_vp_pred,
  output [7:0]  io_master_state_e_1_base_vs1_id,
  output        io_master_state_e_1_base_vs1_valid, io_master_state_e_1_base_vs1_scalar,
  output        io_master_state_e_1_base_vs1_pred,
  output [1:0]  io_master_state_e_1_base_vs1_prec,
  output [7:0]  io_master_state_e_1_base_vs2_id,
  output        io_master_state_e_1_base_vs2_valid, io_master_state_e_1_base_vs2_scalar,
  output        io_master_state_e_1_base_vs2_pred,
  output [1:0]  io_master_state_e_1_base_vs2_prec,
  output [7:0]  io_master_state_e_1_base_vs3_id,
  output        io_master_state_e_1_base_vs3_valid, io_master_state_e_1_base_vs3_scalar,
  output        io_master_state_e_1_base_vs3_pred,
  output [1:0]  io_master_state_e_1_base_vs3_prec,
  output [7:0]  io_master_state_e_1_base_vd_id,
  output        io_master_state_e_1_base_vd_valid, io_master_state_e_1_base_vd_scalar,
  output        io_master_state_e_1_base_vd_pred,
  output [1:0]  io_master_state_e_1_base_vd_prec,
  output        io_master_state_e_1_rate, io_master_state_e_1_active_viu,
  output        io_master_state_e_1_active_vipu, io_master_state_e_1_active_vimu,
  output        io_master_state_e_1_active_vidu, io_master_state_e_1_active_vfmu,
  output        io_master_state_e_1_active_vfdu, io_master_state_e_1_active_vfcu,
  output        io_master_state_e_1_active_vfvu, io_master_state_e_1_active_vrpu,
  output        io_master_state_e_1_active_vrfu, io_master_state_e_1_active_vpu,
  output        io_master_state_e_1_active_vgu, io_master_state_e_1_active_vcu,
  output        io_master_state_e_1_active_vlu, io_master_state_e_1_active_vsu,
  output        io_master_state_e_1_active_vqu, io_master_state_e_1_raw_0,
  output        io_master_state_e_1_raw_1, io_master_state_e_1_raw_2,
  output        io_master_state_e_1_raw_3, io_master_state_e_1_raw_4,
  output        io_master_state_e_1_raw_5, io_master_state_e_1_raw_6,
  output        io_master_state_e_1_raw_7, io_master_state_e_1_war_0,
  output        io_master_state_e_1_war_1, io_master_state_e_1_war_2,
  output        io_master_state_e_1_war_3, io_master_state_e_1_war_4,
  output        io_master_state_e_1_war_5, io_master_state_e_1_war_6,
  output        io_master_state_e_1_war_7, io_master_state_e_1_waw_0,
  output        io_master_state_e_1_waw_1, io_master_state_e_1_waw_2,
  output        io_master_state_e_1_waw_3, io_master_state_e_1_waw_4,
  output        io_master_state_e_1_waw_5, io_master_state_e_1_waw_6,
  output        io_master_state_e_1_waw_7, io_master_state_e_1_last,
  output [1:0]  io_master_state_e_1_rports,
  output [3:0]  io_master_state_e_1_wport_sram,
  output [2:0]  io_master_state_e_1_wport_pred,
  output [9:0]  io_master_state_e_2_fn_union,
  output [63:0] io_master_state_e_2_sreg_ss1, io_master_state_e_2_sreg_ss2,
  output [63:0] io_master_state_e_2_sreg_ss3,
  output [3:0]  io_master_state_e_2_base_vp_id,
  output        io_master_state_e_2_base_vp_valid, io_master_state_e_2_base_vp_scalar,
  output        io_master_state_e_2_base_vp_pred,
  output [7:0]  io_master_state_e_2_base_vs1_id,
  output        io_master_state_e_2_base_vs1_valid, io_master_state_e_2_base_vs1_scalar,
  output        io_master_state_e_2_base_vs1_pred,
  output [1:0]  io_master_state_e_2_base_vs1_prec,
  output [7:0]  io_master_state_e_2_base_vs2_id,
  output        io_master_state_e_2_base_vs2_valid, io_master_state_e_2_base_vs2_scalar,
  output        io_master_state_e_2_base_vs2_pred,
  output [1:0]  io_master_state_e_2_base_vs2_prec,
  output [7:0]  io_master_state_e_2_base_vs3_id,
  output        io_master_state_e_2_base_vs3_valid, io_master_state_e_2_base_vs3_scalar,
  output        io_master_state_e_2_base_vs3_pred,
  output [1:0]  io_master_state_e_2_base_vs3_prec,
  output [7:0]  io_master_state_e_2_base_vd_id,
  output        io_master_state_e_2_base_vd_valid, io_master_state_e_2_base_vd_scalar,
  output        io_master_state_e_2_base_vd_pred,
  output [1:0]  io_master_state_e_2_base_vd_prec,
  output        io_master_state_e_2_rate, io_master_state_e_2_active_viu,
  output        io_master_state_e_2_active_vipu, io_master_state_e_2_active_vimu,
  output        io_master_state_e_2_active_vidu, io_master_state_e_2_active_vfmu,
  output        io_master_state_e_2_active_vfdu, io_master_state_e_2_active_vfcu,
  output        io_master_state_e_2_active_vfvu, io_master_state_e_2_active_vrpu,
  output        io_master_state_e_2_active_vrfu, io_master_state_e_2_active_vpu,
  output        io_master_state_e_2_active_vgu, io_master_state_e_2_active_vcu,
  output        io_master_state_e_2_active_vlu, io_master_state_e_2_active_vsu,
  output        io_master_state_e_2_active_vqu, io_master_state_e_2_raw_0,
  output        io_master_state_e_2_raw_1, io_master_state_e_2_raw_2,
  output        io_master_state_e_2_raw_3, io_master_state_e_2_raw_4,
  output        io_master_state_e_2_raw_5, io_master_state_e_2_raw_6,
  output        io_master_state_e_2_raw_7, io_master_state_e_2_war_0,
  output        io_master_state_e_2_war_1, io_master_state_e_2_war_2,
  output        io_master_state_e_2_war_3, io_master_state_e_2_war_4,
  output        io_master_state_e_2_war_5, io_master_state_e_2_war_6,
  output        io_master_state_e_2_war_7, io_master_state_e_2_waw_0,
  output        io_master_state_e_2_waw_1, io_master_state_e_2_waw_2,
  output        io_master_state_e_2_waw_3, io_master_state_e_2_waw_4,
  output        io_master_state_e_2_waw_5, io_master_state_e_2_waw_6,
  output        io_master_state_e_2_waw_7, io_master_state_e_2_last,
  output [1:0]  io_master_state_e_2_rports,
  output [3:0]  io_master_state_e_2_wport_sram,
  output [2:0]  io_master_state_e_2_wport_pred,
  output [9:0]  io_master_state_e_3_fn_union,
  output [63:0] io_master_state_e_3_sreg_ss1, io_master_state_e_3_sreg_ss2,
  output [63:0] io_master_state_e_3_sreg_ss3,
  output [3:0]  io_master_state_e_3_base_vp_id,
  output        io_master_state_e_3_base_vp_valid, io_master_state_e_3_base_vp_scalar,
  output        io_master_state_e_3_base_vp_pred,
  output [7:0]  io_master_state_e_3_base_vs1_id,
  output        io_master_state_e_3_base_vs1_valid, io_master_state_e_3_base_vs1_scalar,
  output        io_master_state_e_3_base_vs1_pred,
  output [1:0]  io_master_state_e_3_base_vs1_prec,
  output [7:0]  io_master_state_e_3_base_vs2_id,
  output        io_master_state_e_3_base_vs2_valid, io_master_state_e_3_base_vs2_scalar,
  output        io_master_state_e_3_base_vs2_pred,
  output [1:0]  io_master_state_e_3_base_vs2_prec,
  output [7:0]  io_master_state_e_3_base_vs3_id,
  output        io_master_state_e_3_base_vs3_valid, io_master_state_e_3_base_vs3_scalar,
  output        io_master_state_e_3_base_vs3_pred,
  output [1:0]  io_master_state_e_3_base_vs3_prec,
  output [7:0]  io_master_state_e_3_base_vd_id,
  output        io_master_state_e_3_base_vd_valid, io_master_state_e_3_base_vd_scalar,
  output        io_master_state_e_3_base_vd_pred,
  output [1:0]  io_master_state_e_3_base_vd_prec,
  output        io_master_state_e_3_rate, io_master_state_e_3_active_viu,
  output        io_master_state_e_3_active_vipu, io_master_state_e_3_active_vimu,
  output        io_master_state_e_3_active_vidu, io_master_state_e_3_active_vfmu,
  output        io_master_state_e_3_active_vfdu, io_master_state_e_3_active_vfcu,
  output        io_master_state_e_3_active_vfvu, io_master_state_e_3_active_vrpu,
  output        io_master_state_e_3_active_vrfu, io_master_state_e_3_active_vpu,
  output        io_master_state_e_3_active_vgu, io_master_state_e_3_active_vcu,
  output        io_master_state_e_3_active_vlu, io_master_state_e_3_active_vsu,
  output        io_master_state_e_3_active_vqu, io_master_state_e_3_raw_0,
  output        io_master_state_e_3_raw_1, io_master_state_e_3_raw_2,
  output        io_master_state_e_3_raw_3, io_master_state_e_3_raw_4,
  output        io_master_state_e_3_raw_5, io_master_state_e_3_raw_6,
  output        io_master_state_e_3_raw_7, io_master_state_e_3_war_0,
  output        io_master_state_e_3_war_1, io_master_state_e_3_war_2,
  output        io_master_state_e_3_war_3, io_master_state_e_3_war_4,
  output        io_master_state_e_3_war_5, io_master_state_e_3_war_6,
  output        io_master_state_e_3_war_7, io_master_state_e_3_waw_0,
  output        io_master_state_e_3_waw_1, io_master_state_e_3_waw_2,
  output        io_master_state_e_3_waw_3, io_master_state_e_3_waw_4,
  output        io_master_state_e_3_waw_5, io_master_state_e_3_waw_6,
  output        io_master_state_e_3_waw_7, io_master_state_e_3_last,
  output [1:0]  io_master_state_e_3_rports,
  output [3:0]  io_master_state_e_3_wport_sram,
  output [2:0]  io_master_state_e_3_wport_pred,
  output [9:0]  io_master_state_e_4_fn_union,
  output [63:0] io_master_state_e_4_sreg_ss1, io_master_state_e_4_sreg_ss2,
  output [63:0] io_master_state_e_4_sreg_ss3,
  output [3:0]  io_master_state_e_4_base_vp_id,
  output        io_master_state_e_4_base_vp_valid, io_master_state_e_4_base_vp_scalar,
  output        io_master_state_e_4_base_vp_pred,
  output [7:0]  io_master_state_e_4_base_vs1_id,
  output        io_master_state_e_4_base_vs1_valid, io_master_state_e_4_base_vs1_scalar,
  output        io_master_state_e_4_base_vs1_pred,
  output [1:0]  io_master_state_e_4_base_vs1_prec,
  output [7:0]  io_master_state_e_4_base_vs2_id,
  output        io_master_state_e_4_base_vs2_valid, io_master_state_e_4_base_vs2_scalar,
  output        io_master_state_e_4_base_vs2_pred,
  output [1:0]  io_master_state_e_4_base_vs2_prec,
  output [7:0]  io_master_state_e_4_base_vs3_id,
  output        io_master_state_e_4_base_vs3_valid, io_master_state_e_4_base_vs3_scalar,
  output        io_master_state_e_4_base_vs3_pred,
  output [1:0]  io_master_state_e_4_base_vs3_prec,
  output [7:0]  io_master_state_e_4_base_vd_id,
  output        io_master_state_e_4_base_vd_valid, io_master_state_e_4_base_vd_scalar,
  output        io_master_state_e_4_base_vd_pred,
  output [1:0]  io_master_state_e_4_base_vd_prec,
  output        io_master_state_e_4_rate, io_master_state_e_4_active_viu,
  output        io_master_state_e_4_active_vipu, io_master_state_e_4_active_vimu,
  output        io_master_state_e_4_active_vidu, io_master_state_e_4_active_vfmu,
  output        io_master_state_e_4_active_vfdu, io_master_state_e_4_active_vfcu,
  output        io_master_state_e_4_active_vfvu, io_master_state_e_4_active_vrpu,
  output        io_master_state_e_4_active_vrfu, io_master_state_e_4_active_vpu,
  output        io_master_state_e_4_active_vgu, io_master_state_e_4_active_vcu,
  output        io_master_state_e_4_active_vlu, io_master_state_e_4_active_vsu,
  output        io_master_state_e_4_active_vqu, io_master_state_e_4_raw_0,
  output        io_master_state_e_4_raw_1, io_master_state_e_4_raw_2,
  output        io_master_state_e_4_raw_3, io_master_state_e_4_raw_4,
  output        io_master_state_e_4_raw_5, io_master_state_e_4_raw_6,
  output        io_master_state_e_4_raw_7, io_master_state_e_4_war_0,
  output        io_master_state_e_4_war_1, io_master_state_e_4_war_2,
  output        io_master_state_e_4_war_3, io_master_state_e_4_war_4,
  output        io_master_state_e_4_war_5, io_master_state_e_4_war_6,
  output        io_master_state_e_4_war_7, io_master_state_e_4_waw_0,
  output        io_master_state_e_4_waw_1, io_master_state_e_4_waw_2,
  output        io_master_state_e_4_waw_3, io_master_state_e_4_waw_4,
  output        io_master_state_e_4_waw_5, io_master_state_e_4_waw_6,
  output        io_master_state_e_4_waw_7, io_master_state_e_4_last,
  output [1:0]  io_master_state_e_4_rports,
  output [3:0]  io_master_state_e_4_wport_sram,
  output [2:0]  io_master_state_e_4_wport_pred,
  output [9:0]  io_master_state_e_5_fn_union,
  output [63:0] io_master_state_e_5_sreg_ss1, io_master_state_e_5_sreg_ss2,
  output [63:0] io_master_state_e_5_sreg_ss3,
  output [3:0]  io_master_state_e_5_base_vp_id,
  output        io_master_state_e_5_base_vp_valid, io_master_state_e_5_base_vp_scalar,
  output        io_master_state_e_5_base_vp_pred,
  output [7:0]  io_master_state_e_5_base_vs1_id,
  output        io_master_state_e_5_base_vs1_valid, io_master_state_e_5_base_vs1_scalar,
  output        io_master_state_e_5_base_vs1_pred,
  output [1:0]  io_master_state_e_5_base_vs1_prec,
  output [7:0]  io_master_state_e_5_base_vs2_id,
  output        io_master_state_e_5_base_vs2_valid, io_master_state_e_5_base_vs2_scalar,
  output        io_master_state_e_5_base_vs2_pred,
  output [1:0]  io_master_state_e_5_base_vs2_prec,
  output [7:0]  io_master_state_e_5_base_vs3_id,
  output        io_master_state_e_5_base_vs3_valid, io_master_state_e_5_base_vs3_scalar,
  output        io_master_state_e_5_base_vs3_pred,
  output [1:0]  io_master_state_e_5_base_vs3_prec,
  output [7:0]  io_master_state_e_5_base_vd_id,
  output        io_master_state_e_5_base_vd_valid, io_master_state_e_5_base_vd_scalar,
  output        io_master_state_e_5_base_vd_pred,
  output [1:0]  io_master_state_e_5_base_vd_prec,
  output        io_master_state_e_5_rate, io_master_state_e_5_active_viu,
  output        io_master_state_e_5_active_vipu, io_master_state_e_5_active_vimu,
  output        io_master_state_e_5_active_vidu, io_master_state_e_5_active_vfmu,
  output        io_master_state_e_5_active_vfdu, io_master_state_e_5_active_vfcu,
  output        io_master_state_e_5_active_vfvu, io_master_state_e_5_active_vrpu,
  output        io_master_state_e_5_active_vrfu, io_master_state_e_5_active_vpu,
  output        io_master_state_e_5_active_vgu, io_master_state_e_5_active_vcu,
  output        io_master_state_e_5_active_vlu, io_master_state_e_5_active_vsu,
  output        io_master_state_e_5_active_vqu, io_master_state_e_5_raw_0,
  output        io_master_state_e_5_raw_1, io_master_state_e_5_raw_2,
  output        io_master_state_e_5_raw_3, io_master_state_e_5_raw_4,
  output        io_master_state_e_5_raw_5, io_master_state_e_5_raw_6,
  output        io_master_state_e_5_raw_7, io_master_state_e_5_war_0,
  output        io_master_state_e_5_war_1, io_master_state_e_5_war_2,
  output        io_master_state_e_5_war_3, io_master_state_e_5_war_4,
  output        io_master_state_e_5_war_5, io_master_state_e_5_war_6,
  output        io_master_state_e_5_war_7, io_master_state_e_5_waw_0,
  output        io_master_state_e_5_waw_1, io_master_state_e_5_waw_2,
  output        io_master_state_e_5_waw_3, io_master_state_e_5_waw_4,
  output        io_master_state_e_5_waw_5, io_master_state_e_5_waw_6,
  output        io_master_state_e_5_waw_7, io_master_state_e_5_last,
  output [1:0]  io_master_state_e_5_rports,
  output [3:0]  io_master_state_e_5_wport_sram,
  output [2:0]  io_master_state_e_5_wport_pred,
  output [9:0]  io_master_state_e_6_fn_union,
  output [63:0] io_master_state_e_6_sreg_ss1, io_master_state_e_6_sreg_ss2,
  output [63:0] io_master_state_e_6_sreg_ss3,
  output [3:0]  io_master_state_e_6_base_vp_id,
  output        io_master_state_e_6_base_vp_valid, io_master_state_e_6_base_vp_scalar,
  output        io_master_state_e_6_base_vp_pred,
  output [7:0]  io_master_state_e_6_base_vs1_id,
  output        io_master_state_e_6_base_vs1_valid, io_master_state_e_6_base_vs1_scalar,
  output        io_master_state_e_6_base_vs1_pred,
  output [1:0]  io_master_state_e_6_base_vs1_prec,
  output [7:0]  io_master_state_e_6_base_vs2_id,
  output        io_master_state_e_6_base_vs2_valid, io_master_state_e_6_base_vs2_scalar,
  output        io_master_state_e_6_base_vs2_pred,
  output [1:0]  io_master_state_e_6_base_vs2_prec,
  output [7:0]  io_master_state_e_6_base_vs3_id,
  output        io_master_state_e_6_base_vs3_valid, io_master_state_e_6_base_vs3_scalar,
  output        io_master_state_e_6_base_vs3_pred,
  output [1:0]  io_master_state_e_6_base_vs3_prec,
  output [7:0]  io_master_state_e_6_base_vd_id,
  output        io_master_state_e_6_base_vd_valid, io_master_state_e_6_base_vd_scalar,
  output        io_master_state_e_6_base_vd_pred,
  output [1:0]  io_master_state_e_6_base_vd_prec,
  output        io_master_state_e_6_rate, io_master_state_e_6_active_viu,
  output        io_master_state_e_6_active_vipu, io_master_state_e_6_active_vimu,
  output        io_master_state_e_6_active_vidu, io_master_state_e_6_active_vfmu,
  output        io_master_state_e_6_active_vfdu, io_master_state_e_6_active_vfcu,
  output        io_master_state_e_6_active_vfvu, io_master_state_e_6_active_vrpu,
  output        io_master_state_e_6_active_vrfu, io_master_state_e_6_active_vpu,
  output        io_master_state_e_6_active_vgu, io_master_state_e_6_active_vcu,
  output        io_master_state_e_6_active_vlu, io_master_state_e_6_active_vsu,
  output        io_master_state_e_6_active_vqu, io_master_state_e_6_raw_0,
  output        io_master_state_e_6_raw_1, io_master_state_e_6_raw_2,
  output        io_master_state_e_6_raw_3, io_master_state_e_6_raw_4,
  output        io_master_state_e_6_raw_5, io_master_state_e_6_raw_6,
  output        io_master_state_e_6_raw_7, io_master_state_e_6_war_0,
  output        io_master_state_e_6_war_1, io_master_state_e_6_war_2,
  output        io_master_state_e_6_war_3, io_master_state_e_6_war_4,
  output        io_master_state_e_6_war_5, io_master_state_e_6_war_6,
  output        io_master_state_e_6_war_7, io_master_state_e_6_waw_0,
  output        io_master_state_e_6_waw_1, io_master_state_e_6_waw_2,
  output        io_master_state_e_6_waw_3, io_master_state_e_6_waw_4,
  output        io_master_state_e_6_waw_5, io_master_state_e_6_waw_6,
  output        io_master_state_e_6_waw_7, io_master_state_e_6_last,
  output [1:0]  io_master_state_e_6_rports,
  output [3:0]  io_master_state_e_6_wport_sram,
  output [2:0]  io_master_state_e_6_wport_pred,
  output [9:0]  io_master_state_e_7_fn_union,
  output [63:0] io_master_state_e_7_sreg_ss1, io_master_state_e_7_sreg_ss2,
  output [63:0] io_master_state_e_7_sreg_ss3,
  output [3:0]  io_master_state_e_7_base_vp_id,
  output        io_master_state_e_7_base_vp_valid, io_master_state_e_7_base_vp_scalar,
  output        io_master_state_e_7_base_vp_pred,
  output [7:0]  io_master_state_e_7_base_vs1_id,
  output        io_master_state_e_7_base_vs1_valid, io_master_state_e_7_base_vs1_scalar,
  output        io_master_state_e_7_base_vs1_pred,
  output [1:0]  io_master_state_e_7_base_vs1_prec,
  output [7:0]  io_master_state_e_7_base_vs2_id,
  output        io_master_state_e_7_base_vs2_valid, io_master_state_e_7_base_vs2_scalar,
  output        io_master_state_e_7_base_vs2_pred,
  output [1:0]  io_master_state_e_7_base_vs2_prec,
  output [7:0]  io_master_state_e_7_base_vs3_id,
  output        io_master_state_e_7_base_vs3_valid, io_master_state_e_7_base_vs3_scalar,
  output        io_master_state_e_7_base_vs3_pred,
  output [1:0]  io_master_state_e_7_base_vs3_prec,
  output [7:0]  io_master_state_e_7_base_vd_id,
  output        io_master_state_e_7_base_vd_valid, io_master_state_e_7_base_vd_scalar,
  output        io_master_state_e_7_base_vd_pred,
  output [1:0]  io_master_state_e_7_base_vd_prec,
  output        io_master_state_e_7_rate, io_master_state_e_7_active_viu,
  output        io_master_state_e_7_active_vipu, io_master_state_e_7_active_vimu,
  output        io_master_state_e_7_active_vidu, io_master_state_e_7_active_vfmu,
  output        io_master_state_e_7_active_vfdu, io_master_state_e_7_active_vfcu,
  output        io_master_state_e_7_active_vfvu, io_master_state_e_7_active_vrpu,
  output        io_master_state_e_7_active_vrfu, io_master_state_e_7_active_vpu,
  output        io_master_state_e_7_active_vgu, io_master_state_e_7_active_vcu,
  output        io_master_state_e_7_active_vlu, io_master_state_e_7_active_vsu,
  output        io_master_state_e_7_active_vqu, io_master_state_e_7_raw_0,
  output        io_master_state_e_7_raw_1, io_master_state_e_7_raw_2,
  output        io_master_state_e_7_raw_3, io_master_state_e_7_raw_4,
  output        io_master_state_e_7_raw_5, io_master_state_e_7_raw_6,
  output        io_master_state_e_7_raw_7, io_master_state_e_7_war_0,
  output        io_master_state_e_7_war_1, io_master_state_e_7_war_2,
  output        io_master_state_e_7_war_3, io_master_state_e_7_war_4,
  output        io_master_state_e_7_war_5, io_master_state_e_7_war_6,
  output        io_master_state_e_7_war_7, io_master_state_e_7_waw_0,
  output        io_master_state_e_7_waw_1, io_master_state_e_7_waw_2,
  output        io_master_state_e_7_waw_3, io_master_state_e_7_waw_4,
  output        io_master_state_e_7_waw_5, io_master_state_e_7_waw_6,
  output        io_master_state_e_7_waw_7, io_master_state_e_7_last,
  output [1:0]  io_master_state_e_7_rports,
  output [3:0]  io_master_state_e_7_wport_sram,
  output [2:0]  io_master_state_e_7_wport_pred, io_master_state_head,
  output        io_master_update_valid_0, io_master_update_valid_1,
  output        io_master_update_valid_2, io_master_update_valid_3,
  output        io_master_update_valid_4, io_master_update_valid_5,
  output        io_master_update_valid_6, io_master_update_valid_7,
  output [7:0]  io_master_update_reg_0_vp_id, io_master_update_reg_0_vs1_id,
  output [7:0]  io_master_update_reg_0_vs2_id, io_master_update_reg_0_vs3_id,
  output [7:0]  io_master_update_reg_0_vd_id, io_master_update_reg_1_vp_id,
  output [7:0]  io_master_update_reg_1_vs1_id, io_master_update_reg_1_vs2_id,
  output [7:0]  io_master_update_reg_1_vs3_id, io_master_update_reg_1_vd_id,
  output [7:0]  io_master_update_reg_2_vp_id, io_master_update_reg_2_vs1_id,
  output [7:0]  io_master_update_reg_2_vs2_id, io_master_update_reg_2_vs3_id,
  output [7:0]  io_master_update_reg_2_vd_id, io_master_update_reg_3_vp_id,
  output [7:0]  io_master_update_reg_3_vs1_id, io_master_update_reg_3_vs2_id,
  output [7:0]  io_master_update_reg_3_vs3_id, io_master_update_reg_3_vd_id,
  output [7:0]  io_master_update_reg_4_vp_id, io_master_update_reg_4_vs1_id,
  output [7:0]  io_master_update_reg_4_vs2_id, io_master_update_reg_4_vs3_id,
  output [7:0]  io_master_update_reg_4_vd_id, io_master_update_reg_5_vp_id,
  output [7:0]  io_master_update_reg_5_vs1_id, io_master_update_reg_5_vs2_id,
  output [7:0]  io_master_update_reg_5_vs3_id, io_master_update_reg_5_vd_id,
  output [7:0]  io_master_update_reg_6_vp_id, io_master_update_reg_6_vs1_id,
  output [7:0]  io_master_update_reg_6_vs2_id, io_master_update_reg_6_vs3_id,
  output [7:0]  io_master_update_reg_6_vd_id, io_master_update_reg_7_vp_id,
  output [7:0]  io_master_update_reg_7_vs1_id, io_master_update_reg_7_vs2_id,
  output [7:0]  io_master_update_reg_7_vs3_id, io_master_update_reg_7_vd_id,
  output        io_pending_mem, io_pending_all, io_vf_last,
  output [2:0]  io_counters_memoryUOps, io_counters_arithUOps, io_counters_predUOps,
  output [2:0]  io_debug_head, io_debug_tail,
  output        io_debug_maybe_full,
  output [3:0]  io_debug_empty);

  wire        _T;	// sequencer-master.scala:399:66
  reg         casez_tmp;	// sequencer-master.scala:438:21
  reg         casez_tmp_0;	// sequencer-master.scala:438:21
  reg         casez_tmp_1;	// sequencer-master.scala:373:43
  reg         v_0;	// sequencer-master.scala:107:14
  reg         v_1;	// sequencer-master.scala:107:14
  reg         v_2;	// sequencer-master.scala:107:14
  reg         v_3;	// sequencer-master.scala:107:14
  reg         v_4;	// sequencer-master.scala:107:14
  reg         v_5;	// sequencer-master.scala:107:14
  reg         v_6;	// sequencer-master.scala:107:14
  reg         v_7;	// sequencer-master.scala:107:14
  reg  [9:0]  e_0_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_0_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_0_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_0_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_0_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_0_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_0_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_0_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_0_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_0_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_0_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_0_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_0_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_0_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_0_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_0_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_0_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_0_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_0_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_0_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_0_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_0_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_0_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_0_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_0_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_0_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_0_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_0_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_0_active_viu;	// sequencer-master.scala:109:14
  reg         e_0_active_vipu;	// sequencer-master.scala:109:14
  reg         e_0_active_vimu;	// sequencer-master.scala:109:14
  reg         e_0_active_vidu;	// sequencer-master.scala:109:14
  reg         e_0_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_0_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_0_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_0_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_0_active_vpu;	// sequencer-master.scala:109:14
  reg         e_0_active_vgu;	// sequencer-master.scala:109:14
  reg         e_0_active_vcu;	// sequencer-master.scala:109:14
  reg         e_0_active_vlu;	// sequencer-master.scala:109:14
  reg         e_0_active_vsu;	// sequencer-master.scala:109:14
  reg         e_0_active_vqu;	// sequencer-master.scala:109:14
  reg         e_0_raw_0;	// sequencer-master.scala:109:14
  reg         e_0_raw_1;	// sequencer-master.scala:109:14
  reg         e_0_raw_2;	// sequencer-master.scala:109:14
  reg         e_0_raw_3;	// sequencer-master.scala:109:14
  reg         e_0_raw_4;	// sequencer-master.scala:109:14
  reg         e_0_raw_5;	// sequencer-master.scala:109:14
  reg         e_0_raw_6;	// sequencer-master.scala:109:14
  reg         e_0_raw_7;	// sequencer-master.scala:109:14
  reg         e_0_war_0;	// sequencer-master.scala:109:14
  reg         e_0_war_1;	// sequencer-master.scala:109:14
  reg         e_0_war_2;	// sequencer-master.scala:109:14
  reg         e_0_war_3;	// sequencer-master.scala:109:14
  reg         e_0_war_4;	// sequencer-master.scala:109:14
  reg         e_0_war_5;	// sequencer-master.scala:109:14
  reg         e_0_war_6;	// sequencer-master.scala:109:14
  reg         e_0_war_7;	// sequencer-master.scala:109:14
  reg         e_0_waw_0;	// sequencer-master.scala:109:14
  reg         e_0_waw_1;	// sequencer-master.scala:109:14
  reg         e_0_waw_2;	// sequencer-master.scala:109:14
  reg         e_0_waw_3;	// sequencer-master.scala:109:14
  reg         e_0_waw_4;	// sequencer-master.scala:109:14
  reg         e_0_waw_5;	// sequencer-master.scala:109:14
  reg         e_0_waw_6;	// sequencer-master.scala:109:14
  reg         e_0_waw_7;	// sequencer-master.scala:109:14
  reg         e_0_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_0_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_0_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_0_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_1_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_1_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_1_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_1_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_1_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_1_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_1_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_1_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_1_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_1_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_1_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_1_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_1_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_1_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_1_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_1_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_1_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_1_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_1_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_1_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_1_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_1_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_1_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_1_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_1_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_1_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_1_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_1_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_1_active_viu;	// sequencer-master.scala:109:14
  reg         e_1_active_vipu;	// sequencer-master.scala:109:14
  reg         e_1_active_vimu;	// sequencer-master.scala:109:14
  reg         e_1_active_vidu;	// sequencer-master.scala:109:14
  reg         e_1_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_1_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_1_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_1_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_1_active_vpu;	// sequencer-master.scala:109:14
  reg         e_1_active_vgu;	// sequencer-master.scala:109:14
  reg         e_1_active_vcu;	// sequencer-master.scala:109:14
  reg         e_1_active_vlu;	// sequencer-master.scala:109:14
  reg         e_1_active_vsu;	// sequencer-master.scala:109:14
  reg         e_1_active_vqu;	// sequencer-master.scala:109:14
  reg         e_1_raw_0;	// sequencer-master.scala:109:14
  reg         e_1_raw_1;	// sequencer-master.scala:109:14
  reg         e_1_raw_2;	// sequencer-master.scala:109:14
  reg         e_1_raw_3;	// sequencer-master.scala:109:14
  reg         e_1_raw_4;	// sequencer-master.scala:109:14
  reg         e_1_raw_5;	// sequencer-master.scala:109:14
  reg         e_1_raw_6;	// sequencer-master.scala:109:14
  reg         e_1_raw_7;	// sequencer-master.scala:109:14
  reg         e_1_war_0;	// sequencer-master.scala:109:14
  reg         e_1_war_1;	// sequencer-master.scala:109:14
  reg         e_1_war_2;	// sequencer-master.scala:109:14
  reg         e_1_war_3;	// sequencer-master.scala:109:14
  reg         e_1_war_4;	// sequencer-master.scala:109:14
  reg         e_1_war_5;	// sequencer-master.scala:109:14
  reg         e_1_war_6;	// sequencer-master.scala:109:14
  reg         e_1_war_7;	// sequencer-master.scala:109:14
  reg         e_1_waw_0;	// sequencer-master.scala:109:14
  reg         e_1_waw_1;	// sequencer-master.scala:109:14
  reg         e_1_waw_2;	// sequencer-master.scala:109:14
  reg         e_1_waw_3;	// sequencer-master.scala:109:14
  reg         e_1_waw_4;	// sequencer-master.scala:109:14
  reg         e_1_waw_5;	// sequencer-master.scala:109:14
  reg         e_1_waw_6;	// sequencer-master.scala:109:14
  reg         e_1_waw_7;	// sequencer-master.scala:109:14
  reg         e_1_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_1_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_1_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_1_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_2_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_2_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_2_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_2_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_2_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_2_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_2_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_2_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_2_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_2_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_2_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_2_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_2_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_2_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_2_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_2_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_2_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_2_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_2_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_2_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_2_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_2_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_2_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_2_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_2_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_2_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_2_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_2_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_2_active_viu;	// sequencer-master.scala:109:14
  reg         e_2_active_vipu;	// sequencer-master.scala:109:14
  reg         e_2_active_vimu;	// sequencer-master.scala:109:14
  reg         e_2_active_vidu;	// sequencer-master.scala:109:14
  reg         e_2_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_2_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_2_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_2_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_2_active_vpu;	// sequencer-master.scala:109:14
  reg         e_2_active_vgu;	// sequencer-master.scala:109:14
  reg         e_2_active_vcu;	// sequencer-master.scala:109:14
  reg         e_2_active_vlu;	// sequencer-master.scala:109:14
  reg         e_2_active_vsu;	// sequencer-master.scala:109:14
  reg         e_2_active_vqu;	// sequencer-master.scala:109:14
  reg         e_2_raw_0;	// sequencer-master.scala:109:14
  reg         e_2_raw_1;	// sequencer-master.scala:109:14
  reg         e_2_raw_2;	// sequencer-master.scala:109:14
  reg         e_2_raw_3;	// sequencer-master.scala:109:14
  reg         e_2_raw_4;	// sequencer-master.scala:109:14
  reg         e_2_raw_5;	// sequencer-master.scala:109:14
  reg         e_2_raw_6;	// sequencer-master.scala:109:14
  reg         e_2_raw_7;	// sequencer-master.scala:109:14
  reg         e_2_war_0;	// sequencer-master.scala:109:14
  reg         e_2_war_1;	// sequencer-master.scala:109:14
  reg         e_2_war_2;	// sequencer-master.scala:109:14
  reg         e_2_war_3;	// sequencer-master.scala:109:14
  reg         e_2_war_4;	// sequencer-master.scala:109:14
  reg         e_2_war_5;	// sequencer-master.scala:109:14
  reg         e_2_war_6;	// sequencer-master.scala:109:14
  reg         e_2_war_7;	// sequencer-master.scala:109:14
  reg         e_2_waw_0;	// sequencer-master.scala:109:14
  reg         e_2_waw_1;	// sequencer-master.scala:109:14
  reg         e_2_waw_2;	// sequencer-master.scala:109:14
  reg         e_2_waw_3;	// sequencer-master.scala:109:14
  reg         e_2_waw_4;	// sequencer-master.scala:109:14
  reg         e_2_waw_5;	// sequencer-master.scala:109:14
  reg         e_2_waw_6;	// sequencer-master.scala:109:14
  reg         e_2_waw_7;	// sequencer-master.scala:109:14
  reg         e_2_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_2_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_2_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_2_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_3_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_3_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_3_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_3_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_3_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_3_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_3_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_3_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_3_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_3_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_3_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_3_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_3_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_3_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_3_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_3_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_3_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_3_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_3_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_3_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_3_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_3_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_3_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_3_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_3_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_3_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_3_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_3_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_3_active_viu;	// sequencer-master.scala:109:14
  reg         e_3_active_vipu;	// sequencer-master.scala:109:14
  reg         e_3_active_vimu;	// sequencer-master.scala:109:14
  reg         e_3_active_vidu;	// sequencer-master.scala:109:14
  reg         e_3_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_3_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_3_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_3_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_3_active_vpu;	// sequencer-master.scala:109:14
  reg         e_3_active_vgu;	// sequencer-master.scala:109:14
  reg         e_3_active_vcu;	// sequencer-master.scala:109:14
  reg         e_3_active_vlu;	// sequencer-master.scala:109:14
  reg         e_3_active_vsu;	// sequencer-master.scala:109:14
  reg         e_3_active_vqu;	// sequencer-master.scala:109:14
  reg         e_3_raw_0;	// sequencer-master.scala:109:14
  reg         e_3_raw_1;	// sequencer-master.scala:109:14
  reg         e_3_raw_2;	// sequencer-master.scala:109:14
  reg         e_3_raw_3;	// sequencer-master.scala:109:14
  reg         e_3_raw_4;	// sequencer-master.scala:109:14
  reg         e_3_raw_5;	// sequencer-master.scala:109:14
  reg         e_3_raw_6;	// sequencer-master.scala:109:14
  reg         e_3_raw_7;	// sequencer-master.scala:109:14
  reg         e_3_war_0;	// sequencer-master.scala:109:14
  reg         e_3_war_1;	// sequencer-master.scala:109:14
  reg         e_3_war_2;	// sequencer-master.scala:109:14
  reg         e_3_war_3;	// sequencer-master.scala:109:14
  reg         e_3_war_4;	// sequencer-master.scala:109:14
  reg         e_3_war_5;	// sequencer-master.scala:109:14
  reg         e_3_war_6;	// sequencer-master.scala:109:14
  reg         e_3_war_7;	// sequencer-master.scala:109:14
  reg         e_3_waw_0;	// sequencer-master.scala:109:14
  reg         e_3_waw_1;	// sequencer-master.scala:109:14
  reg         e_3_waw_2;	// sequencer-master.scala:109:14
  reg         e_3_waw_3;	// sequencer-master.scala:109:14
  reg         e_3_waw_4;	// sequencer-master.scala:109:14
  reg         e_3_waw_5;	// sequencer-master.scala:109:14
  reg         e_3_waw_6;	// sequencer-master.scala:109:14
  reg         e_3_waw_7;	// sequencer-master.scala:109:14
  reg         e_3_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_3_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_3_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_3_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_4_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_4_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_4_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_4_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_4_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_4_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_4_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_4_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_4_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_4_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_4_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_4_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_4_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_4_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_4_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_4_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_4_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_4_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_4_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_4_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_4_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_4_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_4_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_4_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_4_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_4_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_4_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_4_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_4_active_viu;	// sequencer-master.scala:109:14
  reg         e_4_active_vipu;	// sequencer-master.scala:109:14
  reg         e_4_active_vimu;	// sequencer-master.scala:109:14
  reg         e_4_active_vidu;	// sequencer-master.scala:109:14
  reg         e_4_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_4_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_4_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_4_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_4_active_vpu;	// sequencer-master.scala:109:14
  reg         e_4_active_vgu;	// sequencer-master.scala:109:14
  reg         e_4_active_vcu;	// sequencer-master.scala:109:14
  reg         e_4_active_vlu;	// sequencer-master.scala:109:14
  reg         e_4_active_vsu;	// sequencer-master.scala:109:14
  reg         e_4_active_vqu;	// sequencer-master.scala:109:14
  reg         e_4_raw_0;	// sequencer-master.scala:109:14
  reg         e_4_raw_1;	// sequencer-master.scala:109:14
  reg         e_4_raw_2;	// sequencer-master.scala:109:14
  reg         e_4_raw_3;	// sequencer-master.scala:109:14
  reg         e_4_raw_4;	// sequencer-master.scala:109:14
  reg         e_4_raw_5;	// sequencer-master.scala:109:14
  reg         e_4_raw_6;	// sequencer-master.scala:109:14
  reg         e_4_raw_7;	// sequencer-master.scala:109:14
  reg         e_4_war_0;	// sequencer-master.scala:109:14
  reg         e_4_war_1;	// sequencer-master.scala:109:14
  reg         e_4_war_2;	// sequencer-master.scala:109:14
  reg         e_4_war_3;	// sequencer-master.scala:109:14
  reg         e_4_war_4;	// sequencer-master.scala:109:14
  reg         e_4_war_5;	// sequencer-master.scala:109:14
  reg         e_4_war_6;	// sequencer-master.scala:109:14
  reg         e_4_war_7;	// sequencer-master.scala:109:14
  reg         e_4_waw_0;	// sequencer-master.scala:109:14
  reg         e_4_waw_1;	// sequencer-master.scala:109:14
  reg         e_4_waw_2;	// sequencer-master.scala:109:14
  reg         e_4_waw_3;	// sequencer-master.scala:109:14
  reg         e_4_waw_4;	// sequencer-master.scala:109:14
  reg         e_4_waw_5;	// sequencer-master.scala:109:14
  reg         e_4_waw_6;	// sequencer-master.scala:109:14
  reg         e_4_waw_7;	// sequencer-master.scala:109:14
  reg         e_4_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_4_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_4_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_4_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_5_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_5_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_5_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_5_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_5_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_5_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_5_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_5_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_5_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_5_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_5_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_5_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_5_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_5_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_5_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_5_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_5_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_5_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_5_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_5_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_5_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_5_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_5_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_5_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_5_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_5_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_5_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_5_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_5_active_viu;	// sequencer-master.scala:109:14
  reg         e_5_active_vipu;	// sequencer-master.scala:109:14
  reg         e_5_active_vimu;	// sequencer-master.scala:109:14
  reg         e_5_active_vidu;	// sequencer-master.scala:109:14
  reg         e_5_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_5_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_5_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_5_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_5_active_vpu;	// sequencer-master.scala:109:14
  reg         e_5_active_vgu;	// sequencer-master.scala:109:14
  reg         e_5_active_vcu;	// sequencer-master.scala:109:14
  reg         e_5_active_vlu;	// sequencer-master.scala:109:14
  reg         e_5_active_vsu;	// sequencer-master.scala:109:14
  reg         e_5_active_vqu;	// sequencer-master.scala:109:14
  reg         e_5_raw_0;	// sequencer-master.scala:109:14
  reg         e_5_raw_1;	// sequencer-master.scala:109:14
  reg         e_5_raw_2;	// sequencer-master.scala:109:14
  reg         e_5_raw_3;	// sequencer-master.scala:109:14
  reg         e_5_raw_4;	// sequencer-master.scala:109:14
  reg         e_5_raw_5;	// sequencer-master.scala:109:14
  reg         e_5_raw_6;	// sequencer-master.scala:109:14
  reg         e_5_raw_7;	// sequencer-master.scala:109:14
  reg         e_5_war_0;	// sequencer-master.scala:109:14
  reg         e_5_war_1;	// sequencer-master.scala:109:14
  reg         e_5_war_2;	// sequencer-master.scala:109:14
  reg         e_5_war_3;	// sequencer-master.scala:109:14
  reg         e_5_war_4;	// sequencer-master.scala:109:14
  reg         e_5_war_5;	// sequencer-master.scala:109:14
  reg         e_5_war_6;	// sequencer-master.scala:109:14
  reg         e_5_war_7;	// sequencer-master.scala:109:14
  reg         e_5_waw_0;	// sequencer-master.scala:109:14
  reg         e_5_waw_1;	// sequencer-master.scala:109:14
  reg         e_5_waw_2;	// sequencer-master.scala:109:14
  reg         e_5_waw_3;	// sequencer-master.scala:109:14
  reg         e_5_waw_4;	// sequencer-master.scala:109:14
  reg         e_5_waw_5;	// sequencer-master.scala:109:14
  reg         e_5_waw_6;	// sequencer-master.scala:109:14
  reg         e_5_waw_7;	// sequencer-master.scala:109:14
  reg         e_5_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_5_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_5_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_5_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_6_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_6_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_6_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_6_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_6_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_6_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_6_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_6_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_6_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_6_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_6_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_6_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_6_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_6_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_6_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_6_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_6_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_6_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_6_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_6_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_6_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_6_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_6_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_6_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_6_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_6_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_6_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_6_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_6_active_viu;	// sequencer-master.scala:109:14
  reg         e_6_active_vipu;	// sequencer-master.scala:109:14
  reg         e_6_active_vimu;	// sequencer-master.scala:109:14
  reg         e_6_active_vidu;	// sequencer-master.scala:109:14
  reg         e_6_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_6_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_6_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_6_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_6_active_vpu;	// sequencer-master.scala:109:14
  reg         e_6_active_vgu;	// sequencer-master.scala:109:14
  reg         e_6_active_vcu;	// sequencer-master.scala:109:14
  reg         e_6_active_vlu;	// sequencer-master.scala:109:14
  reg         e_6_active_vsu;	// sequencer-master.scala:109:14
  reg         e_6_active_vqu;	// sequencer-master.scala:109:14
  reg         e_6_raw_0;	// sequencer-master.scala:109:14
  reg         e_6_raw_1;	// sequencer-master.scala:109:14
  reg         e_6_raw_2;	// sequencer-master.scala:109:14
  reg         e_6_raw_3;	// sequencer-master.scala:109:14
  reg         e_6_raw_4;	// sequencer-master.scala:109:14
  reg         e_6_raw_5;	// sequencer-master.scala:109:14
  reg         e_6_raw_6;	// sequencer-master.scala:109:14
  reg         e_6_raw_7;	// sequencer-master.scala:109:14
  reg         e_6_war_0;	// sequencer-master.scala:109:14
  reg         e_6_war_1;	// sequencer-master.scala:109:14
  reg         e_6_war_2;	// sequencer-master.scala:109:14
  reg         e_6_war_3;	// sequencer-master.scala:109:14
  reg         e_6_war_4;	// sequencer-master.scala:109:14
  reg         e_6_war_5;	// sequencer-master.scala:109:14
  reg         e_6_war_6;	// sequencer-master.scala:109:14
  reg         e_6_war_7;	// sequencer-master.scala:109:14
  reg         e_6_waw_0;	// sequencer-master.scala:109:14
  reg         e_6_waw_1;	// sequencer-master.scala:109:14
  reg         e_6_waw_2;	// sequencer-master.scala:109:14
  reg         e_6_waw_3;	// sequencer-master.scala:109:14
  reg         e_6_waw_4;	// sequencer-master.scala:109:14
  reg         e_6_waw_5;	// sequencer-master.scala:109:14
  reg         e_6_waw_6;	// sequencer-master.scala:109:14
  reg         e_6_waw_7;	// sequencer-master.scala:109:14
  reg         e_6_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_6_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_6_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_6_wport_pred;	// sequencer-master.scala:109:14
  reg  [9:0]  e_7_fn_union;	// sequencer-master.scala:109:14
  reg  [63:0] e_7_sreg_ss1;	// sequencer-master.scala:109:14
  reg  [63:0] e_7_sreg_ss2;	// sequencer-master.scala:109:14
  reg  [63:0] e_7_sreg_ss3;	// sequencer-master.scala:109:14
  reg  [3:0]  e_7_base_vp_id;	// sequencer-master.scala:109:14
  reg         e_7_base_vp_valid;	// sequencer-master.scala:109:14
  reg         e_7_base_vp_scalar;	// sequencer-master.scala:109:14
  reg         e_7_base_vp_pred;	// sequencer-master.scala:109:14
  reg  [7:0]  e_7_base_vs1_id;	// sequencer-master.scala:109:14
  reg         e_7_base_vs1_valid;	// sequencer-master.scala:109:14
  reg         e_7_base_vs1_scalar;	// sequencer-master.scala:109:14
  reg         e_7_base_vs1_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_7_base_vs1_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_7_base_vs2_id;	// sequencer-master.scala:109:14
  reg         e_7_base_vs2_valid;	// sequencer-master.scala:109:14
  reg         e_7_base_vs2_scalar;	// sequencer-master.scala:109:14
  reg         e_7_base_vs2_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_7_base_vs2_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_7_base_vs3_id;	// sequencer-master.scala:109:14
  reg         e_7_base_vs3_valid;	// sequencer-master.scala:109:14
  reg         e_7_base_vs3_scalar;	// sequencer-master.scala:109:14
  reg         e_7_base_vs3_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_7_base_vs3_prec;	// sequencer-master.scala:109:14
  reg  [7:0]  e_7_base_vd_id;	// sequencer-master.scala:109:14
  reg         e_7_base_vd_valid;	// sequencer-master.scala:109:14
  reg         e_7_base_vd_scalar;	// sequencer-master.scala:109:14
  reg         e_7_base_vd_pred;	// sequencer-master.scala:109:14
  reg  [1:0]  e_7_base_vd_prec;	// sequencer-master.scala:109:14
  reg         e_7_active_viu;	// sequencer-master.scala:109:14
  reg         e_7_active_vipu;	// sequencer-master.scala:109:14
  reg         e_7_active_vimu;	// sequencer-master.scala:109:14
  reg         e_7_active_vidu;	// sequencer-master.scala:109:14
  reg         e_7_active_vfmu;	// sequencer-master.scala:109:14
  reg         e_7_active_vfdu;	// sequencer-master.scala:109:14
  reg         e_7_active_vfcu;	// sequencer-master.scala:109:14
  reg         e_7_active_vfvu;	// sequencer-master.scala:109:14
  reg         e_7_active_vpu;	// sequencer-master.scala:109:14
  reg         e_7_active_vgu;	// sequencer-master.scala:109:14
  reg         e_7_active_vcu;	// sequencer-master.scala:109:14
  reg         e_7_active_vlu;	// sequencer-master.scala:109:14
  reg         e_7_active_vsu;	// sequencer-master.scala:109:14
  reg         e_7_active_vqu;	// sequencer-master.scala:109:14
  reg         e_7_raw_0;	// sequencer-master.scala:109:14
  reg         e_7_raw_1;	// sequencer-master.scala:109:14
  reg         e_7_raw_2;	// sequencer-master.scala:109:14
  reg         e_7_raw_3;	// sequencer-master.scala:109:14
  reg         e_7_raw_4;	// sequencer-master.scala:109:14
  reg         e_7_raw_5;	// sequencer-master.scala:109:14
  reg         e_7_raw_6;	// sequencer-master.scala:109:14
  reg         e_7_raw_7;	// sequencer-master.scala:109:14
  reg         e_7_war_0;	// sequencer-master.scala:109:14
  reg         e_7_war_1;	// sequencer-master.scala:109:14
  reg         e_7_war_2;	// sequencer-master.scala:109:14
  reg         e_7_war_3;	// sequencer-master.scala:109:14
  reg         e_7_war_4;	// sequencer-master.scala:109:14
  reg         e_7_war_5;	// sequencer-master.scala:109:14
  reg         e_7_war_6;	// sequencer-master.scala:109:14
  reg         e_7_war_7;	// sequencer-master.scala:109:14
  reg         e_7_waw_0;	// sequencer-master.scala:109:14
  reg         e_7_waw_1;	// sequencer-master.scala:109:14
  reg         e_7_waw_2;	// sequencer-master.scala:109:14
  reg         e_7_waw_3;	// sequencer-master.scala:109:14
  reg         e_7_waw_4;	// sequencer-master.scala:109:14
  reg         e_7_waw_5;	// sequencer-master.scala:109:14
  reg         e_7_waw_6;	// sequencer-master.scala:109:14
  reg         e_7_waw_7;	// sequencer-master.scala:109:14
  reg         e_7_last;	// sequencer-master.scala:109:14
  reg  [1:0]  e_7_rports;	// sequencer-master.scala:109:14
  reg  [3:0]  e_7_wport_sram;	// sequencer-master.scala:109:14
  reg  [2:0]  e_7_wport_pred;	// sequencer-master.scala:109:14
  reg         maybe_full;	// sequencer-master.scala:111:23
  reg  [2:0]  head;	// sequencer-master.scala:112:17
  reg  [2:0]  tail;	// sequencer-master.scala:113:17
  reg         _T_2_398;	// sequencer-master.scala:444:24

  wire [2:0] _T_0 = tail + 3'h1;	// sequencer-master.scala:267:35, util.scala:94:11
  wire [2:0] _T_1 = tail + 3'h2;	// sequencer-master.scala:267:35, util.scala:94:11
  wire [2:0] _T_2 = tail + 3'h3;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_3 = _T & io_op_valid;	// Decoupled.scala:37:37, sequencer-master.scala:399:66
  wire _T_4 = tail == 3'h0;	// sequencer-master.scala:112:17, :267:35, util.scala:94:11
  wire _T_5 = tail == 3'h1;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_6 = tail == 3'h2;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_7 = tail == 3'h3;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_8 = tail == 3'h4;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_9 = tail == 3'h5;	// sequencer-master.scala:183:52, :267:35, util.scala:94:11
  wire _T_10 = tail == 3'h6;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_11 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire _T_12 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire _T_13 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire _T_14 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire _T_15 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire _T_16 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire _T_17 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire _T_18 = io_op_bits_active_vint & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire _T_19 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_20 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_21 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_22 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_23 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_24 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_25 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_26 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_27 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_28 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_29 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_30 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_31 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_32 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_33 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_34 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_35 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:364:41
  wire _T_36 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:364:41
  wire _T_37 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:364:41
  wire _T_38 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:364:41
  wire _T_39 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:364:41
  wire _T_40 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:364:41
  wire _T_41 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:364:41
  wire _T_42 = io_op_bits_active_vint & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :364:41, util.scala:94:11
  wire [7:0] _T_43 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_4 | _T_19 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_19 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_44 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_5 | _T_20 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_20 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_45 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_6 | _T_21 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_21 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_46 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_7 | _T_22 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_22 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_47 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_8 | _T_23 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_23 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_48 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_9 | _T_24 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_24 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_49 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_10 | _T_25 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_25 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_50 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (&tail | _T_26 ?
                io_op_bits_reg_vs1_id : 8'h0) : _T_26 ? io_op_bits_reg_vs1_id : 8'h0;	// sequencer-master.scala:267:35, :330:47, :411:70, util.scala:94:11
  wire [7:0] _T_51 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_4 | _T_27 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_27 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_52 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_5 | _T_28 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_28 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_53 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_6 | _T_29 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_29 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_54 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_7 | _T_30 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_30 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_55 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_8 | _T_31 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_31 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_56 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_9 | _T_32 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_32 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_57 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_10 | _T_33 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_33 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:330:47, :411:70
  wire [7:0] _T_58 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (&tail | _T_34 ?
                io_op_bits_reg_vs2_id : 8'h0) : _T_34 ? io_op_bits_reg_vs2_id : 8'h0;	// sequencer-master.scala:267:35, :330:47, :411:70, util.scala:94:11
  wire _T_59 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_60 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_61 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_62 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_63 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_64 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_65 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_66 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_67 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_4 | _T_35 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_35 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_68 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_5 | _T_36 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_36 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_69 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_6 | _T_37 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_37 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_70 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_7 | _T_38 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_38 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_71 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_8 | _T_39 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_39 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_72 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_9 | _T_40 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_40 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_73 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_10 | _T_41 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_41 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:364:41, :411:70
  wire [7:0] _T_74 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (&tail | _T_42 ? io_op_bits_reg_vd_id
                : 8'h0) : _T_42 ? io_op_bits_reg_vd_id : 8'h0;	// sequencer-master.scala:267:35, :364:41, :411:70, util.scala:94:11
  wire [7:0] _T_75 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_4 | _T_11 ? io_op_bits_reg_vp_id :
                8'h0) : _T_11 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_76 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_5 | _T_12 ? io_op_bits_reg_vp_id :
                8'h0) : _T_12 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_77 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_6 | _T_13 ? io_op_bits_reg_vp_id :
                8'h0) : _T_13 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_78 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_7 | _T_14 ? io_op_bits_reg_vp_id :
                8'h0) : _T_14 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_79 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_8 | _T_15 ? io_op_bits_reg_vp_id :
                8'h0) : _T_15 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_80 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_9 | _T_16 ? io_op_bits_reg_vp_id :
                8'h0) : _T_16 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_81 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_10 | _T_17 ? io_op_bits_reg_vp_id
                : 8'h0) : _T_17 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:322:41, :411:70
  wire [7:0] _T_82 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (&tail | _T_18 ? io_op_bits_reg_vp_id
                : 8'h0) : _T_18 ? io_op_bits_reg_vp_id : 8'h0;	// sequencer-master.scala:267:35, :322:41, :411:70, util.scala:94:11
  wire _T_83 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_84 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_85 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_86 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_87 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_88 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_89 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_90 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_91 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_92 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_93 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_94 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_95 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_96 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_97 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_98 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_99 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:364:41
  wire _T_100 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:364:41
  wire _T_101 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:364:41
  wire _T_102 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:364:41
  wire _T_103 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:364:41
  wire _T_104 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:364:41
  wire _T_105 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:364:41
  wire _T_106 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :364:41, util.scala:94:11
  wire _T_107 = io_op_bits_active_vidiv | io_op_bits_active_vfdiv;	// sequencer-master.scala:298:31
  wire _T_108 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire _T_109 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire _T_110 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire _T_111 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire _T_112 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire _T_113 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire _T_114 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire _T_115 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_116 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_83 ? io_op_bits_reg_vs1_id
                : _T_43) : _T_83 ? io_op_bits_reg_vs1_id : _T_43;	// sequencer-master.scala:330:47
  wire [7:0] _T_117 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_84 ? io_op_bits_reg_vs1_id
                : _T_44) : _T_84 ? io_op_bits_reg_vs1_id : _T_44;	// sequencer-master.scala:330:47
  wire [7:0] _T_118 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_85 ? io_op_bits_reg_vs1_id
                : _T_45) : _T_85 ? io_op_bits_reg_vs1_id : _T_45;	// sequencer-master.scala:330:47
  wire [7:0] _T_119 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_86 ? io_op_bits_reg_vs1_id
                : _T_46) : _T_86 ? io_op_bits_reg_vs1_id : _T_46;	// sequencer-master.scala:330:47
  wire [7:0] _T_120 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_87 ? io_op_bits_reg_vs1_id
                : _T_47) : _T_87 ? io_op_bits_reg_vs1_id : _T_47;	// sequencer-master.scala:330:47
  wire [7:0] _T_121 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_88 ? io_op_bits_reg_vs1_id
                : _T_48) : _T_88 ? io_op_bits_reg_vs1_id : _T_48;	// sequencer-master.scala:330:47
  wire [7:0] _T_122 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_89 ?
                io_op_bits_reg_vs1_id : _T_49) : _T_89 ? io_op_bits_reg_vs1_id : _T_49;	// sequencer-master.scala:330:47
  wire [7:0] _T_123 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (&tail | _T_90 ?
                io_op_bits_reg_vs1_id : _T_50) : _T_90 ? io_op_bits_reg_vs1_id : _T_50;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_124 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_91 ? io_op_bits_reg_vs2_id
                : _T_51) : _T_91 ? io_op_bits_reg_vs2_id : _T_51;	// sequencer-master.scala:330:47
  wire [7:0] _T_125 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_92 ? io_op_bits_reg_vs2_id
                : _T_52) : _T_92 ? io_op_bits_reg_vs2_id : _T_52;	// sequencer-master.scala:330:47
  wire [7:0] _T_126 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_93 ? io_op_bits_reg_vs2_id
                : _T_53) : _T_93 ? io_op_bits_reg_vs2_id : _T_53;	// sequencer-master.scala:330:47
  wire [7:0] _T_127 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_94 ? io_op_bits_reg_vs2_id
                : _T_54) : _T_94 ? io_op_bits_reg_vs2_id : _T_54;	// sequencer-master.scala:330:47
  wire [7:0] _T_128 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_95 ? io_op_bits_reg_vs2_id
                : _T_55) : _T_95 ? io_op_bits_reg_vs2_id : _T_55;	// sequencer-master.scala:330:47
  wire [7:0] _T_129 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_96 ? io_op_bits_reg_vs2_id
                : _T_56) : _T_96 ? io_op_bits_reg_vs2_id : _T_56;	// sequencer-master.scala:330:47
  wire [7:0] _T_130 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_97 ?
                io_op_bits_reg_vs2_id : _T_57) : _T_97 ? io_op_bits_reg_vs2_id : _T_57;	// sequencer-master.scala:330:47
  wire [7:0] _T_131 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (&tail | _T_98 ?
                io_op_bits_reg_vs2_id : _T_58) : _T_98 ? io_op_bits_reg_vs2_id : _T_58;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_132 = _T_0 == 3'h0;	// sequencer-master.scala:112:17, :267:35
  wire _T_133 = _T_0 == 3'h1;	// sequencer-master.scala:267:35
  wire _T_134 = _T_0 == 3'h2;	// sequencer-master.scala:267:35
  wire _T_135 = _T_0 == 3'h3;	// sequencer-master.scala:267:35
  wire _T_136 = _T_0 == 3'h4;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_137 = _T_0 == 3'h5;	// sequencer-master.scala:183:52, :267:35
  wire _T_138 = _T_0 == 3'h6;	// sequencer-master.scala:267:35
  wire [7:0] _T_139 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_132 | _T_99 ? io_op_bits_reg_vd_id
                : _T_67) : _T_99 ? io_op_bits_reg_vd_id : _T_67;	// sequencer-master.scala:364:41
  wire [7:0] _T_140 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_133 | _T_100 ?
                io_op_bits_reg_vd_id : _T_68) : _T_100 ? io_op_bits_reg_vd_id : _T_68;	// sequencer-master.scala:364:41
  wire [7:0] _T_141 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_134 | _T_101 ?
                io_op_bits_reg_vd_id : _T_69) : _T_101 ? io_op_bits_reg_vd_id : _T_69;	// sequencer-master.scala:364:41
  wire [7:0] _T_142 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_135 | _T_102 ?
                io_op_bits_reg_vd_id : _T_70) : _T_102 ? io_op_bits_reg_vd_id : _T_70;	// sequencer-master.scala:364:41
  wire [7:0] _T_143 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_136 | _T_103 ?
                io_op_bits_reg_vd_id : _T_71) : _T_103 ? io_op_bits_reg_vd_id : _T_71;	// sequencer-master.scala:364:41
  wire [7:0] _T_144 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_137 | _T_104 ?
                io_op_bits_reg_vd_id : _T_72) : _T_104 ? io_op_bits_reg_vd_id : _T_72;	// sequencer-master.scala:364:41
  wire [7:0] _T_145 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_138 | _T_105 ?
                io_op_bits_reg_vd_id : _T_73) : _T_105 ? io_op_bits_reg_vd_id : _T_73;	// sequencer-master.scala:364:41
  wire [7:0] _T_146 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_106 ? io_op_bits_reg_vd_id
                : _T_74) : _T_106 ? io_op_bits_reg_vd_id : _T_74;	// sequencer-master.scala:267:35, :364:41
  wire [7:0] _T_147 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_4 | _T_108 ? io_op_bits_reg_vp_id :
                _T_75) : _T_108 ? io_op_bits_reg_vp_id : _T_75;	// sequencer-master.scala:322:41
  wire [7:0] _T_148 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_5 | _T_109 ? io_op_bits_reg_vp_id :
                _T_76) : _T_109 ? io_op_bits_reg_vp_id : _T_76;	// sequencer-master.scala:322:41
  wire [7:0] _T_149 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_6 | _T_110 ? io_op_bits_reg_vp_id :
                _T_77) : _T_110 ? io_op_bits_reg_vp_id : _T_77;	// sequencer-master.scala:322:41
  wire [7:0] _T_150 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_7 | _T_111 ? io_op_bits_reg_vp_id :
                _T_78) : _T_111 ? io_op_bits_reg_vp_id : _T_78;	// sequencer-master.scala:322:41
  wire [7:0] _T_151 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_8 | _T_112 ? io_op_bits_reg_vp_id :
                _T_79) : _T_112 ? io_op_bits_reg_vp_id : _T_79;	// sequencer-master.scala:322:41
  wire [7:0] _T_152 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_9 | _T_113 ? io_op_bits_reg_vp_id :
                _T_80) : _T_113 ? io_op_bits_reg_vp_id : _T_80;	// sequencer-master.scala:322:41
  wire [7:0] _T_153 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_10 | _T_114 ? io_op_bits_reg_vp_id
                : _T_81) : _T_114 ? io_op_bits_reg_vp_id : _T_81;	// sequencer-master.scala:322:41
  wire [7:0] _T_154 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (&tail | _T_115 ? io_op_bits_reg_vp_id
                : _T_82) : _T_115 ? io_op_bits_reg_vp_id : _T_82;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire _T_155 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_156 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_157 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_158 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_159 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_160 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_161 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_162 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_163 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_164 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_165 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_166 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_167 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_168 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_169 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_170 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_171 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:364:41
  wire _T_172 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:364:41
  wire _T_173 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:364:41
  wire _T_174 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:364:41
  wire _T_175 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:364:41
  wire _T_176 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:364:41
  wire _T_177 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:364:41
  wire _T_178 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :364:41, util.scala:94:11
  wire _T_179 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire _T_180 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire _T_181 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire _T_182 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire _T_183 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire _T_184 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire _T_185 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire _T_186 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_187 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_155 ?
                io_op_bits_reg_vs1_id : _T_116) : _T_155 ? io_op_bits_reg_vs1_id : _T_116;	// sequencer-master.scala:330:47
  wire [7:0] _T_188 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_156 ?
                io_op_bits_reg_vs1_id : _T_117) : _T_156 ? io_op_bits_reg_vs1_id : _T_117;	// sequencer-master.scala:330:47
  wire [7:0] _T_189 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_157 ?
                io_op_bits_reg_vs1_id : _T_118) : _T_157 ? io_op_bits_reg_vs1_id : _T_118;	// sequencer-master.scala:330:47
  wire [7:0] _T_190 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_158 ?
                io_op_bits_reg_vs1_id : _T_119) : _T_158 ? io_op_bits_reg_vs1_id : _T_119;	// sequencer-master.scala:330:47
  wire [7:0] _T_191 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_159 ?
                io_op_bits_reg_vs1_id : _T_120) : _T_159 ? io_op_bits_reg_vs1_id : _T_120;	// sequencer-master.scala:330:47
  wire [7:0] _T_192 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_160 ?
                io_op_bits_reg_vs1_id : _T_121) : _T_160 ? io_op_bits_reg_vs1_id : _T_121;	// sequencer-master.scala:330:47
  wire [7:0] _T_193 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_161 ?
                io_op_bits_reg_vs1_id : _T_122) : _T_161 ? io_op_bits_reg_vs1_id : _T_122;	// sequencer-master.scala:330:47
  wire [7:0] _T_194 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (&tail | _T_162 ?
                io_op_bits_reg_vs1_id : _T_123) : _T_162 ? io_op_bits_reg_vs1_id : _T_123;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_195 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_132 | _T_171 ?
                io_op_bits_reg_vd_id : _T_139) : _T_171 ? io_op_bits_reg_vd_id : _T_139;	// sequencer-master.scala:364:41
  wire [7:0] _T_196 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_133 | _T_172 ?
                io_op_bits_reg_vd_id : _T_140) : _T_172 ? io_op_bits_reg_vd_id : _T_140;	// sequencer-master.scala:364:41
  wire [7:0] _T_197 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_134 | _T_173 ?
                io_op_bits_reg_vd_id : _T_141) : _T_173 ? io_op_bits_reg_vd_id : _T_141;	// sequencer-master.scala:364:41
  wire [7:0] _T_198 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_135 | _T_174 ?
                io_op_bits_reg_vd_id : _T_142) : _T_174 ? io_op_bits_reg_vd_id : _T_142;	// sequencer-master.scala:364:41
  wire [7:0] _T_199 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_136 | _T_175 ?
                io_op_bits_reg_vd_id : _T_143) : _T_175 ? io_op_bits_reg_vd_id : _T_143;	// sequencer-master.scala:364:41
  wire [7:0] _T_200 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_137 | _T_176 ?
                io_op_bits_reg_vd_id : _T_144) : _T_176 ? io_op_bits_reg_vd_id : _T_144;	// sequencer-master.scala:364:41
  wire [7:0] _T_201 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_138 | _T_177 ?
                io_op_bits_reg_vd_id : _T_145) : _T_177 ? io_op_bits_reg_vd_id : _T_145;	// sequencer-master.scala:364:41
  wire [7:0] _T_202 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_178 ? io_op_bits_reg_vd_id
                : _T_146) : _T_178 ? io_op_bits_reg_vd_id : _T_146;	// sequencer-master.scala:267:35, :364:41
  wire [7:0] _T_203 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_4 | _T_179 ? io_op_bits_reg_vp_id
                : _T_147) : _T_179 ? io_op_bits_reg_vp_id : _T_147;	// sequencer-master.scala:322:41
  wire [7:0] _T_204 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_5 | _T_180 ? io_op_bits_reg_vp_id
                : _T_148) : _T_180 ? io_op_bits_reg_vp_id : _T_148;	// sequencer-master.scala:322:41
  wire [7:0] _T_205 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_6 | _T_181 ? io_op_bits_reg_vp_id
                : _T_149) : _T_181 ? io_op_bits_reg_vp_id : _T_149;	// sequencer-master.scala:322:41
  wire [7:0] _T_206 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_7 | _T_182 ? io_op_bits_reg_vp_id
                : _T_150) : _T_182 ? io_op_bits_reg_vp_id : _T_150;	// sequencer-master.scala:322:41
  wire [7:0] _T_207 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_8 | _T_183 ? io_op_bits_reg_vp_id
                : _T_151) : _T_183 ? io_op_bits_reg_vp_id : _T_151;	// sequencer-master.scala:322:41
  wire [7:0] _T_208 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_9 | _T_184 ? io_op_bits_reg_vp_id
                : _T_152) : _T_184 ? io_op_bits_reg_vp_id : _T_152;	// sequencer-master.scala:322:41
  wire [7:0] _T_209 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_10 | _T_185 ? io_op_bits_reg_vp_id
                : _T_153) : _T_185 ? io_op_bits_reg_vp_id : _T_153;	// sequencer-master.scala:322:41
  wire [7:0] _T_210 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (&tail | _T_186 ? io_op_bits_reg_vp_id
                : _T_154) : _T_186 ? io_op_bits_reg_vp_id : _T_154;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire _T_211 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:330:47
  wire _T_212 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:330:47
  wire _T_213 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:330:47
  wire _T_214 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:330:47
  wire _T_215 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:330:47
  wire _T_216 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:330:47
  wire _T_217 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:330:47
  wire _T_218 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_219 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:364:41
  wire _T_220 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:364:41
  wire _T_221 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:364:41
  wire _T_222 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:364:41
  wire _T_223 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:364:41
  wire _T_224 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:364:41
  wire _T_225 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:364:41
  wire _T_226 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :364:41, util.scala:94:11
  wire _T_227 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire _T_228 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire _T_229 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire _T_230 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire _T_231 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire _T_232 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire _T_233 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire _T_234 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_235 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_4 | _T_211 ?
                io_op_bits_reg_vs1_id : _T_187) : _T_211 ? io_op_bits_reg_vs1_id : _T_187;	// sequencer-master.scala:330:47
  wire [7:0] _T_236 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_5 | _T_212 ?
                io_op_bits_reg_vs1_id : _T_188) : _T_212 ? io_op_bits_reg_vs1_id : _T_188;	// sequencer-master.scala:330:47
  wire [7:0] _T_237 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_6 | _T_213 ?
                io_op_bits_reg_vs1_id : _T_189) : _T_213 ? io_op_bits_reg_vs1_id : _T_189;	// sequencer-master.scala:330:47
  wire [7:0] _T_238 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_7 | _T_214 ?
                io_op_bits_reg_vs1_id : _T_190) : _T_214 ? io_op_bits_reg_vs1_id : _T_190;	// sequencer-master.scala:330:47
  wire [7:0] _T_239 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_8 | _T_215 ?
                io_op_bits_reg_vs1_id : _T_191) : _T_215 ? io_op_bits_reg_vs1_id : _T_191;	// sequencer-master.scala:330:47
  wire [7:0] _T_240 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_9 | _T_216 ?
                io_op_bits_reg_vs1_id : _T_192) : _T_216 ? io_op_bits_reg_vs1_id : _T_192;	// sequencer-master.scala:330:47
  wire [7:0] _T_241 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_10 | _T_217 ?
                io_op_bits_reg_vs1_id : _T_193) : _T_217 ? io_op_bits_reg_vs1_id : _T_193;	// sequencer-master.scala:330:47
  wire [7:0] _T_242 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (&tail | _T_218 ?
                io_op_bits_reg_vs1_id : _T_194) : _T_218 ? io_op_bits_reg_vs1_id : _T_194;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_243 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_4 | _T_219 ? io_op_bits_reg_vd_id
                : _T_195) : _T_219 ? io_op_bits_reg_vd_id : _T_195;	// sequencer-master.scala:364:41
  wire [7:0] _T_244 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_5 | _T_220 ? io_op_bits_reg_vd_id
                : _T_196) : _T_220 ? io_op_bits_reg_vd_id : _T_196;	// sequencer-master.scala:364:41
  wire [7:0] _T_245 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_6 | _T_221 ? io_op_bits_reg_vd_id
                : _T_197) : _T_221 ? io_op_bits_reg_vd_id : _T_197;	// sequencer-master.scala:364:41
  wire [7:0] _T_246 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_7 | _T_222 ? io_op_bits_reg_vd_id
                : _T_198) : _T_222 ? io_op_bits_reg_vd_id : _T_198;	// sequencer-master.scala:364:41
  wire [7:0] _T_247 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_8 | _T_223 ? io_op_bits_reg_vd_id
                : _T_199) : _T_223 ? io_op_bits_reg_vd_id : _T_199;	// sequencer-master.scala:364:41
  wire [7:0] _T_248 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_9 | _T_224 ? io_op_bits_reg_vd_id
                : _T_200) : _T_224 ? io_op_bits_reg_vd_id : _T_200;	// sequencer-master.scala:364:41
  wire [7:0] _T_249 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_10 | _T_225 ?
                io_op_bits_reg_vd_id : _T_201) : _T_225 ? io_op_bits_reg_vd_id : _T_201;	// sequencer-master.scala:364:41
  wire [7:0] _T_250 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (&tail | _T_226 ?
                io_op_bits_reg_vd_id : _T_202) : _T_226 ? io_op_bits_reg_vd_id : _T_202;	// sequencer-master.scala:267:35, :364:41, util.scala:94:11
  wire [7:0] _T_251 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_4 | _T_227 ? io_op_bits_reg_vp_id
                : _T_203) : _T_227 ? io_op_bits_reg_vp_id : _T_203;	// sequencer-master.scala:322:41
  wire [7:0] _T_252 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_5 | _T_228 ? io_op_bits_reg_vp_id
                : _T_204) : _T_228 ? io_op_bits_reg_vp_id : _T_204;	// sequencer-master.scala:322:41
  wire [7:0] _T_253 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_6 | _T_229 ? io_op_bits_reg_vp_id
                : _T_205) : _T_229 ? io_op_bits_reg_vp_id : _T_205;	// sequencer-master.scala:322:41
  wire [7:0] _T_254 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_7 | _T_230 ? io_op_bits_reg_vp_id
                : _T_206) : _T_230 ? io_op_bits_reg_vp_id : _T_206;	// sequencer-master.scala:322:41
  wire [7:0] _T_255 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_8 | _T_231 ? io_op_bits_reg_vp_id
                : _T_207) : _T_231 ? io_op_bits_reg_vp_id : _T_207;	// sequencer-master.scala:322:41
  wire [7:0] _T_256 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_9 | _T_232 ? io_op_bits_reg_vp_id
                : _T_208) : _T_232 ? io_op_bits_reg_vp_id : _T_208;	// sequencer-master.scala:322:41
  wire [7:0] _T_257 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_10 | _T_233 ?
                io_op_bits_reg_vp_id : _T_209) : _T_233 ? io_op_bits_reg_vp_id : _T_209;	// sequencer-master.scala:322:41
  wire [7:0] _T_258 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (&tail | _T_234 ?
                io_op_bits_reg_vp_id : _T_210) : _T_234 ? io_op_bits_reg_vp_id : _T_210;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire _T_259 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire [7:0] _T_260 = _T_259 ? io_op_bits_reg_vp_id : _T_251;	// sequencer-master.scala:322:41
  wire _T_261 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire [7:0] _T_262 = _T_261 ? io_op_bits_reg_vp_id : _T_252;	// sequencer-master.scala:322:41
  wire _T_263 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire [7:0] _T_264 = _T_263 ? io_op_bits_reg_vp_id : _T_253;	// sequencer-master.scala:322:41
  wire _T_265 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire [7:0] _T_266 = _T_265 ? io_op_bits_reg_vp_id : _T_254;	// sequencer-master.scala:322:41
  wire _T_267 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire [7:0] _T_268 = _T_267 ? io_op_bits_reg_vp_id : _T_255;	// sequencer-master.scala:322:41
  wire _T_269 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire [7:0] _T_270 = _T_269 ? io_op_bits_reg_vp_id : _T_256;	// sequencer-master.scala:322:41
  wire _T_271 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire [7:0] _T_272 = _T_271 ? io_op_bits_reg_vp_id : _T_257;	// sequencer-master.scala:322:41
  wire _T_273 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_274 = _T_273 ? io_op_bits_reg_vp_id : _T_258;	// sequencer-master.scala:322:41
  wire _T_275 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:330:47
  wire [7:0] _T_276 = _T_275 ? io_op_bits_reg_vs1_id : _T_235;	// sequencer-master.scala:330:47
  wire _T_277 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:330:47
  wire [7:0] _T_278 = _T_277 ? io_op_bits_reg_vs1_id : _T_236;	// sequencer-master.scala:330:47
  wire _T_279 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:330:47
  wire [7:0] _T_280 = _T_279 ? io_op_bits_reg_vs1_id : _T_237;	// sequencer-master.scala:330:47
  wire _T_281 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:330:47
  wire [7:0] _T_282 = _T_281 ? io_op_bits_reg_vs1_id : _T_238;	// sequencer-master.scala:330:47
  wire _T_283 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:330:47
  wire [7:0] _T_284 = _T_283 ? io_op_bits_reg_vs1_id : _T_239;	// sequencer-master.scala:330:47
  wire _T_285 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:330:47
  wire [7:0] _T_286 = _T_285 ? io_op_bits_reg_vs1_id : _T_240;	// sequencer-master.scala:330:47
  wire _T_287 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:330:47
  wire [7:0] _T_288 = _T_287 ? io_op_bits_reg_vs1_id : _T_241;	// sequencer-master.scala:330:47
  wire _T_289 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_290 = _T_289 ? io_op_bits_reg_vs1_id : _T_242;	// sequencer-master.scala:330:47
  wire _T_291 = _T_1 == 3'h0;	// sequencer-master.scala:112:17, :267:35
  wire _T_292 = _T_1 == 3'h1;	// sequencer-master.scala:267:35
  wire _T_293 = _T_1 == 3'h2;	// sequencer-master.scala:267:35
  wire _T_294 = _T_1 == 3'h3;	// sequencer-master.scala:267:35
  wire _T_295 = _T_1 == 3'h4;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_296 = _T_1 == 3'h5;	// sequencer-master.scala:183:52, :267:35
  wire _T_297 = _T_1 == 3'h6;	// sequencer-master.scala:267:35
  wire [7:0] _T_298 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_4 | _T_259 ? io_op_bits_reg_vp_id : _T_251) : _T_260) :
                _T_260;	// sequencer-master.scala:322:41
  wire [7:0] _T_299 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_5 | _T_261 ? io_op_bits_reg_vp_id : _T_252) : _T_262) :
                _T_262;	// sequencer-master.scala:322:41
  wire [7:0] _T_300 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_6 | _T_263 ? io_op_bits_reg_vp_id : _T_253) : _T_264) :
                _T_264;	// sequencer-master.scala:322:41
  wire [7:0] _T_301 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_7 | _T_265 ? io_op_bits_reg_vp_id : _T_254) : _T_266) :
                _T_266;	// sequencer-master.scala:322:41
  wire [7:0] _T_302 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_8 | _T_267 ? io_op_bits_reg_vp_id : _T_255) : _T_268) :
                _T_268;	// sequencer-master.scala:322:41
  wire [7:0] _T_303 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_9 | _T_269 ? io_op_bits_reg_vp_id : _T_256) : _T_270) :
                _T_270;	// sequencer-master.scala:322:41
  wire [7:0] _T_304 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_10 | _T_271 ? io_op_bits_reg_vp_id : _T_257) : _T_272) :
                _T_272;	// sequencer-master.scala:322:41
  wire [7:0] _T_305 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (&tail | _T_273 ? io_op_bits_reg_vp_id : _T_258) : _T_274) :
                _T_274;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_306 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_291 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_4 | _T_275 ? io_op_bits_reg_vs1_id : _T_235) : _T_276) :
                _T_276;	// sequencer-master.scala:330:47
  wire [7:0] _T_307 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_292 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_5 | _T_277 ? io_op_bits_reg_vs1_id : _T_236) : _T_278) :
                _T_278;	// sequencer-master.scala:330:47
  wire [7:0] _T_308 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_293 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_6 | _T_279 ? io_op_bits_reg_vs1_id : _T_237) : _T_280) :
                _T_280;	// sequencer-master.scala:330:47
  wire [7:0] _T_309 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_294 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_7 | _T_281 ? io_op_bits_reg_vs1_id : _T_238) : _T_282) :
                _T_282;	// sequencer-master.scala:330:47
  wire [7:0] _T_310 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_295 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_8 | _T_283 ? io_op_bits_reg_vs1_id : _T_239) : _T_284) :
                _T_284;	// sequencer-master.scala:330:47
  wire [7:0] _T_311 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_296 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_9 | _T_285 ? io_op_bits_reg_vs1_id : _T_240) : _T_286) :
                _T_286;	// sequencer-master.scala:330:47
  wire [7:0] _T_312 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_297 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_10 | _T_287 ? io_op_bits_reg_vs1_id : _T_241) : _T_288) :
                _T_288;	// sequencer-master.scala:330:47
  wire [7:0] _T_313 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & &_T_1 ? io_op_bits_reg_vs2_id :
                io_op_bits_base_vs1_valid ? (&tail | _T_289 ? io_op_bits_reg_vs1_id : _T_242) : _T_290) :
                _T_290;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire _T_314 = _T_2 == 3'h0;	// sequencer-master.scala:112:17, :267:35
  wire _T_315 = _T_2 == 3'h1;	// sequencer-master.scala:267:35
  wire _T_316 = _T_2 == 3'h2;	// sequencer-master.scala:267:35
  wire _T_317 = _T_2 == 3'h3;	// sequencer-master.scala:267:35
  wire _T_318 = _T_2 == 3'h4;	// sequencer-master.scala:267:35, util.scala:94:11
  wire _T_319 = _T_2 == 3'h5;	// sequencer-master.scala:183:52, :267:35
  wire _T_320 = _T_2 == 3'h6;	// sequencer-master.scala:267:35
  wire _T_321 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_314;	// sequencer-master.scala:364:41
  wire _T_322 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_315;	// sequencer-master.scala:364:41
  wire _T_323 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_316;	// sequencer-master.scala:364:41
  wire _T_324 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_317;	// sequencer-master.scala:364:41
  wire _T_325 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_318;	// sequencer-master.scala:364:41
  wire _T_326 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_319;	// sequencer-master.scala:364:41
  wire _T_327 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_320;	// sequencer-master.scala:364:41
  wire _T_328 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & &_T_2;	// sequencer-master.scala:267:35, :364:41
  wire _T_329 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire [7:0] _T_330 = _T_329 ? io_op_bits_reg_vp_id : _T_298;	// sequencer-master.scala:322:41
  wire _T_331 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire [7:0] _T_332 = _T_331 ? io_op_bits_reg_vp_id : _T_299;	// sequencer-master.scala:322:41
  wire _T_333 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire [7:0] _T_334 = _T_333 ? io_op_bits_reg_vp_id : _T_300;	// sequencer-master.scala:322:41
  wire _T_335 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire [7:0] _T_336 = _T_335 ? io_op_bits_reg_vp_id : _T_301;	// sequencer-master.scala:322:41
  wire _T_337 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire [7:0] _T_338 = _T_337 ? io_op_bits_reg_vp_id : _T_302;	// sequencer-master.scala:322:41
  wire _T_339 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire [7:0] _T_340 = _T_339 ? io_op_bits_reg_vp_id : _T_303;	// sequencer-master.scala:322:41
  wire _T_341 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire [7:0] _T_342 = _T_341 ? io_op_bits_reg_vp_id : _T_304;	// sequencer-master.scala:322:41
  wire _T_343 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_344 = _T_343 ? io_op_bits_reg_vp_id : _T_305;	// sequencer-master.scala:322:41
  wire _T_345 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:330:47
  wire [7:0] _T_346 = _T_345 ? io_op_bits_reg_vs2_id : _T_306;	// sequencer-master.scala:330:47
  wire _T_347 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:330:47
  wire [7:0] _T_348 = _T_347 ? io_op_bits_reg_vs2_id : _T_307;	// sequencer-master.scala:330:47
  wire _T_349 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:330:47
  wire [7:0] _T_350 = _T_349 ? io_op_bits_reg_vs2_id : _T_308;	// sequencer-master.scala:330:47
  wire _T_351 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:330:47
  wire [7:0] _T_352 = _T_351 ? io_op_bits_reg_vs2_id : _T_309;	// sequencer-master.scala:330:47
  wire _T_353 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:330:47
  wire [7:0] _T_354 = _T_353 ? io_op_bits_reg_vs2_id : _T_310;	// sequencer-master.scala:330:47
  wire _T_355 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:330:47
  wire [7:0] _T_356 = _T_355 ? io_op_bits_reg_vs2_id : _T_311;	// sequencer-master.scala:330:47
  wire _T_357 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:330:47
  wire [7:0] _T_358 = _T_357 ? io_op_bits_reg_vs2_id : _T_312;	// sequencer-master.scala:330:47
  wire _T_359 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :330:47, util.scala:94:11
  wire [7:0] _T_360 = _T_359 ? io_op_bits_reg_vs2_id : _T_313;	// sequencer-master.scala:330:47
  wire [7:0] _T_361 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_4 | _T_329 ? io_op_bits_reg_vp_id : _T_298) : _T_330) :
                _T_330;	// sequencer-master.scala:322:41
  wire [7:0] _T_362 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_5 | _T_331 ? io_op_bits_reg_vp_id : _T_299) : _T_332) :
                _T_332;	// sequencer-master.scala:322:41
  wire [7:0] _T_363 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_6 | _T_333 ? io_op_bits_reg_vp_id : _T_300) : _T_334) :
                _T_334;	// sequencer-master.scala:322:41
  wire [7:0] _T_364 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_7 | _T_335 ? io_op_bits_reg_vp_id : _T_301) : _T_336) :
                _T_336;	// sequencer-master.scala:322:41
  wire [7:0] _T_365 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_8 | _T_337 ? io_op_bits_reg_vp_id : _T_302) : _T_338) :
                _T_338;	// sequencer-master.scala:322:41
  wire [7:0] _T_366 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_9 | _T_339 ? io_op_bits_reg_vp_id : _T_303) : _T_340) :
                _T_340;	// sequencer-master.scala:322:41
  wire [7:0] _T_367 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_10 | _T_341 ? io_op_bits_reg_vp_id : _T_304) : _T_342) :
                _T_342;	// sequencer-master.scala:322:41
  wire [7:0] _T_368 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (&tail | _T_343 ? io_op_bits_reg_vp_id : _T_305) : _T_344) :
                _T_344;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire _T_369 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:322:41
  wire [7:0] _T_370 = _T_369 ? io_op_bits_reg_vp_id : _T_361;	// sequencer-master.scala:322:41
  wire _T_371 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:322:41
  wire [7:0] _T_372 = _T_371 ? io_op_bits_reg_vp_id : _T_362;	// sequencer-master.scala:322:41
  wire _T_373 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:322:41
  wire [7:0] _T_374 = _T_373 ? io_op_bits_reg_vp_id : _T_363;	// sequencer-master.scala:322:41
  wire _T_375 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:322:41
  wire [7:0] _T_376 = _T_375 ? io_op_bits_reg_vp_id : _T_364;	// sequencer-master.scala:322:41
  wire _T_377 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:322:41
  wire [7:0] _T_378 = _T_377 ? io_op_bits_reg_vp_id : _T_365;	// sequencer-master.scala:322:41
  wire _T_379 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:322:41
  wire [7:0] _T_380 = _T_379 ? io_op_bits_reg_vp_id : _T_366;	// sequencer-master.scala:322:41
  wire _T_381 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:322:41
  wire [7:0] _T_382 = _T_381 ? io_op_bits_reg_vp_id : _T_367;	// sequencer-master.scala:322:41
  wire _T_383 = io_op_bits_active_vld & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :322:41, util.scala:94:11
  wire [7:0] _T_384 = _T_383 ? io_op_bits_reg_vp_id : _T_368;	// sequencer-master.scala:322:41
  wire _T_385 = _T_3 & (io_op_bits_active_vst & (_T_291 | _T_132 | _T_4) | io_op_bits_active_vld & (_T_291
                | _T_132 | _T_4) | io_op_bits_active_vstx & (_T_291 | _T_132 | _T_4) |
                io_op_bits_active_vldx & (_T_291 | _T_132 | _T_4) | io_op_bits_active_vamo & (_T_314 |
                _T_291 | _T_132 | _T_4) | io_op_bits_active_vrfirst & _T_4 | io_op_bits_active_vrpred &
                _T_4 | io_op_bits_active_vfconv & _T_4 | io_op_bits_active_vfcmp & _T_4 |
                io_op_bits_active_vfdiv & (_T_132 | _T_4) | io_op_bits_active_vfma & _T_4 |
                io_op_bits_active_vidiv & (_T_132 | _T_4) | io_op_bits_active_vimul & _T_4 |
                io_op_bits_active_vipred & _T_4 | io_op_bits_active_vint & _T_4);	// sequencer-master.scala:188:42
  wire _T_386 = _T_3 & (io_op_bits_active_vst & (_T_292 | _T_133 | _T_5) | io_op_bits_active_vld & (_T_292
                | _T_133 | _T_5) | io_op_bits_active_vstx & (_T_292 | _T_133 | _T_5) |
                io_op_bits_active_vldx & (_T_292 | _T_133 | _T_5) | io_op_bits_active_vamo & (_T_315 |
                _T_292 | _T_133 | _T_5) | io_op_bits_active_vrfirst & _T_5 | io_op_bits_active_vrpred &
                _T_5 | io_op_bits_active_vfconv & _T_5 | io_op_bits_active_vfcmp & _T_5 |
                io_op_bits_active_vfdiv & (_T_133 | _T_5) | io_op_bits_active_vfma & _T_5 |
                io_op_bits_active_vidiv & (_T_133 | _T_5) | io_op_bits_active_vimul & _T_5 |
                io_op_bits_active_vipred & _T_5 | io_op_bits_active_vint & _T_5);	// sequencer-master.scala:188:42
  wire _T_387 = _T_3 & (io_op_bits_active_vst & (_T_293 | _T_134 | _T_6) | io_op_bits_active_vld & (_T_293
                | _T_134 | _T_6) | io_op_bits_active_vstx & (_T_293 | _T_134 | _T_6) |
                io_op_bits_active_vldx & (_T_293 | _T_134 | _T_6) | io_op_bits_active_vamo & (_T_316 |
                _T_293 | _T_134 | _T_6) | io_op_bits_active_vrfirst & _T_6 | io_op_bits_active_vrpred &
                _T_6 | io_op_bits_active_vfconv & _T_6 | io_op_bits_active_vfcmp & _T_6 |
                io_op_bits_active_vfdiv & (_T_134 | _T_6) | io_op_bits_active_vfma & _T_6 |
                io_op_bits_active_vidiv & (_T_134 | _T_6) | io_op_bits_active_vimul & _T_6 |
                io_op_bits_active_vipred & _T_6 | io_op_bits_active_vint & _T_6);	// sequencer-master.scala:188:42
  wire _T_388 = _T_3 & (io_op_bits_active_vst & (_T_294 | _T_135 | _T_7) | io_op_bits_active_vld & (_T_294
                | _T_135 | _T_7) | io_op_bits_active_vstx & (_T_294 | _T_135 | _T_7) |
                io_op_bits_active_vldx & (_T_294 | _T_135 | _T_7) | io_op_bits_active_vamo & (_T_317 |
                _T_294 | _T_135 | _T_7) | io_op_bits_active_vrfirst & _T_7 | io_op_bits_active_vrpred &
                _T_7 | io_op_bits_active_vfconv & _T_7 | io_op_bits_active_vfcmp & _T_7 |
                io_op_bits_active_vfdiv & (_T_135 | _T_7) | io_op_bits_active_vfma & _T_7 |
                io_op_bits_active_vidiv & (_T_135 | _T_7) | io_op_bits_active_vimul & _T_7 |
                io_op_bits_active_vipred & _T_7 | io_op_bits_active_vint & _T_7);	// sequencer-master.scala:188:42
  wire _T_389 = _T_3 & (io_op_bits_active_vst & (_T_295 | _T_136 | _T_8) | io_op_bits_active_vld & (_T_295
                | _T_136 | _T_8) | io_op_bits_active_vstx & (_T_295 | _T_136 | _T_8) |
                io_op_bits_active_vldx & (_T_295 | _T_136 | _T_8) | io_op_bits_active_vamo & (_T_318 |
                _T_295 | _T_136 | _T_8) | io_op_bits_active_vrfirst & _T_8 | io_op_bits_active_vrpred &
                _T_8 | io_op_bits_active_vfconv & _T_8 | io_op_bits_active_vfcmp & _T_8 |
                io_op_bits_active_vfdiv & (_T_136 | _T_8) | io_op_bits_active_vfma & _T_8 |
                io_op_bits_active_vidiv & (_T_136 | _T_8) | io_op_bits_active_vimul & _T_8 |
                io_op_bits_active_vipred & _T_8 | io_op_bits_active_vint & _T_8);	// sequencer-master.scala:188:42
  wire _T_390 = _T_3 & (io_op_bits_active_vst & (_T_296 | _T_137 | _T_9) | io_op_bits_active_vld & (_T_296
                | _T_137 | _T_9) | io_op_bits_active_vstx & (_T_296 | _T_137 | _T_9) |
                io_op_bits_active_vldx & (_T_296 | _T_137 | _T_9) | io_op_bits_active_vamo & (_T_319 |
                _T_296 | _T_137 | _T_9) | io_op_bits_active_vrfirst & _T_9 | io_op_bits_active_vrpred &
                _T_9 | io_op_bits_active_vfconv & _T_9 | io_op_bits_active_vfcmp & _T_9 |
                io_op_bits_active_vfdiv & (_T_137 | _T_9) | io_op_bits_active_vfma & _T_9 |
                io_op_bits_active_vidiv & (_T_137 | _T_9) | io_op_bits_active_vimul & _T_9 |
                io_op_bits_active_vipred & _T_9 | io_op_bits_active_vint & _T_9);	// sequencer-master.scala:188:42
  wire _T_391 = _T_3 & (io_op_bits_active_vst & (_T_297 | _T_138 | _T_10) | io_op_bits_active_vld & (_T_297
                | _T_138 | _T_10) | io_op_bits_active_vstx & (_T_297 | _T_138 | _T_10) |
                io_op_bits_active_vldx & (_T_297 | _T_138 | _T_10) | io_op_bits_active_vamo & (_T_320 |
                _T_297 | _T_138 | _T_10) | io_op_bits_active_vrfirst & _T_10 | io_op_bits_active_vrpred &
                _T_10 | io_op_bits_active_vfconv & _T_10 | io_op_bits_active_vfcmp & _T_10 |
                io_op_bits_active_vfdiv & (_T_138 | _T_10) | io_op_bits_active_vfma & _T_10 |
                io_op_bits_active_vidiv & (_T_138 | _T_10) | io_op_bits_active_vimul & _T_10 |
                io_op_bits_active_vipred & _T_10 | io_op_bits_active_vint & _T_10);	// sequencer-master.scala:188:42
  wire _T_392 = _T_3 & (io_op_bits_active_vst & (&_T_1 | &_T_0 | &tail) | io_op_bits_active_vld & (&_T_1 |
                &_T_0 | &tail) | io_op_bits_active_vstx & (&_T_1 | &_T_0 | &tail) | io_op_bits_active_vldx
                & (&_T_1 | &_T_0 | &tail) | io_op_bits_active_vamo & (&_T_2 | &_T_1 | &_T_0 | &tail) |
                io_op_bits_active_vrfirst & &tail | io_op_bits_active_vrpred & &tail |
                io_op_bits_active_vfconv & &tail | io_op_bits_active_vfcmp & &tail |
                io_op_bits_active_vfdiv & (&_T_0 | &tail) | io_op_bits_active_vfma & &tail |
                io_op_bits_active_vidiv & (&_T_0 | &tail) | io_op_bits_active_vimul & &tail |
                io_op_bits_active_vipred & &tail | io_op_bits_active_vint & &tail);	// sequencer-master.scala:188:42, :267:35, util.scala:94:11
  wire _T_393 = ~maybe_full & head == tail;	// sequencer-master.scala:389:{15,27,36}, util.scala:94:11
  wire [2:0] _T_394 = head - tail;	// sequencer-master.scala:389:{36,52}, util.scala:94:11
  wire [3:0] _T_395 = {_T_393, _T_394};	// Cat.scala:30:58
  assign _T = |_T_395 & (io_op_bits_active_vint | io_op_bits_active_vipred | io_op_bits_active_vimul |
                io_op_bits_active_vfma | io_op_bits_active_vfcmp | io_op_bits_active_vfconv |
                io_op_bits_active_vrpred | io_op_bits_active_vrfirst) | |{_T_393, _T_394[2:1]} & _T_107 |
                _T_395 > 4'h2 & (io_op_bits_active_vld | io_op_bits_active_vst | io_op_bits_active_vldx |
                io_op_bits_active_vstx) | |{_T_393, _T_394[2]} & io_op_bits_active_vamo;	// sequencer-master.scala:397:{14,26,105}, :398:{14,26}, :399:{14,26,55,66}, :400:{14,26}, util.scala:94:11
  wire [2:0] _T_396 = head + 3'h1;	// sequencer-master.scala:267:35, :389:36, util.scala:94:11
  always @(*) begin	// sequencer-master.scala:438:21
    casez (head)	// sequencer-master.scala:389:36, :438:21
      3'b000:
        casez_tmp = v_0;	// sequencer-master.scala:136:44, :438:21
      3'b001:
        casez_tmp = v_1;	// sequencer-master.scala:136:44, :438:21
      3'b010:
        casez_tmp = v_2;	// sequencer-master.scala:136:44, :438:21
      3'b011:
        casez_tmp = v_3;	// sequencer-master.scala:136:44, :438:21
      3'b100:
        casez_tmp = v_4;	// sequencer-master.scala:136:44, :438:21
      3'b101:
        casez_tmp = v_5;	// sequencer-master.scala:136:44, :438:21
      3'b110:
        casez_tmp = v_6;	// sequencer-master.scala:136:44, :438:21
      default:
        casez_tmp = v_7;	// sequencer-master.scala:136:44, :438:21
    endcase	// sequencer-master.scala:389:36, :438:21
  end // always @(*)
  always @(*) begin	// sequencer-master.scala:438:21
    casez (head)	// sequencer-master.scala:389:36, :438:21
      3'b000:
        casez_tmp_0 = io_master_clear_0;	// sequencer-master.scala:438:21
      3'b001:
        casez_tmp_0 = io_master_clear_1;	// sequencer-master.scala:438:21
      3'b010:
        casez_tmp_0 = io_master_clear_2;	// sequencer-master.scala:438:21
      3'b011:
        casez_tmp_0 = io_master_clear_3;	// sequencer-master.scala:438:21
      3'b100:
        casez_tmp_0 = io_master_clear_4;	// sequencer-master.scala:438:21
      3'b101:
        casez_tmp_0 = io_master_clear_5;	// sequencer-master.scala:438:21
      3'b110:
        casez_tmp_0 = io_master_clear_6;	// sequencer-master.scala:438:21
      default:
        casez_tmp_0 = io_master_clear_7;	// sequencer-master.scala:438:21
    endcase	// sequencer-master.scala:389:36, :438:21
  end // always @(*)
  wire _T_397 = casez_tmp & casez_tmp_0;	// sequencer-master.scala:438:21
  always @(*) begin	// sequencer-master.scala:373:43, :438:21
    casez (head)	// sequencer-master.scala:373:43, :389:36, :438:21
      3'b000:
        casez_tmp_1 = e_0_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b001:
        casez_tmp_1 = e_1_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b010:
        casez_tmp_1 = e_2_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b011:
        casez_tmp_1 = e_3_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b100:
        casez_tmp_1 = e_4_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b101:
        casez_tmp_1 = e_5_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      3'b110:
        casez_tmp_1 = e_6_last;	// sequencer-master.scala:283:19, :373:43, :438:21
      default:
        casez_tmp_1 = e_7_last;	// sequencer-master.scala:283:19, :373:43, :438:21
    endcase	// sequencer-master.scala:373:43, :389:36, :438:21
  end // always @(*)
  `ifndef SYNTHESIS	// sequencer-master.scala:107:14
    `ifdef RANDOMIZE_REG_INIT	// sequencer-master.scala:107:14
      reg [31:0] _RANDOM;	// sequencer-master.scala:107:14
      reg [31:0] _RANDOM_3;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_4;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_5;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_6;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_7;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_8;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_9;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_10;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_11;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_12;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_13;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_14;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_15;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_16;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_17;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_18;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_19;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_20;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_21;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_22;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_23;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_24;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_25;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_26;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_27;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_28;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_29;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_30;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_31;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_32;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_33;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_34;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_35;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_36;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_37;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_38;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_39;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_40;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_41;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_42;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_43;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_44;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_45;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_46;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_47;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_48;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_49;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_50;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_51;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_52;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_53;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_54;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_55;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_56;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_57;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_58;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_59;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_60;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_61;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_62;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_63;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_64;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_65;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_66;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_67;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_68;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_69;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_70;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_71;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_72;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_73;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_74;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_75;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_76;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_77;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_78;	// sequencer-master.scala:109:14
      reg [31:0] _RANDOM_79;	// sequencer-master.scala:109:14

    `endif
    initial begin	// sequencer-master.scala:107:14
      `INIT_RANDOM_PROLOG_	// sequencer-master.scala:107:14
      `ifdef RANDOMIZE_REG_INIT	// sequencer-master.scala:107:14
        _RANDOM = `RANDOM;	// sequencer-master.scala:107:14
        v_0 = _RANDOM[0];	// sequencer-master.scala:107:14
        v_1 = _RANDOM[1];	// sequencer-master.scala:107:14
        v_2 = _RANDOM[2];	// sequencer-master.scala:107:14
        v_3 = _RANDOM[3];	// sequencer-master.scala:107:14
        v_4 = _RANDOM[4];	// sequencer-master.scala:107:14
        v_5 = _RANDOM[5];	// sequencer-master.scala:107:14
        v_6 = _RANDOM[6];	// sequencer-master.scala:107:14
        v_7 = _RANDOM[7];	// sequencer-master.scala:107:14
        e_0_fn_union = _RANDOM[17:8];	// sequencer-master.scala:109:14
        _RANDOM_3 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_4 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_sreg_ss1 = {_RANDOM_4[17:0], _RANDOM_3, _RANDOM[31:18]};	// sequencer-master.scala:109:14
        _RANDOM_5 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_6 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_sreg_ss2 = {_RANDOM_6[17:0], _RANDOM_5, _RANDOM_4[31:18]};	// sequencer-master.scala:109:14
        _RANDOM_7 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_8 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_sreg_ss3 = {_RANDOM_8[17:0], _RANDOM_7, _RANDOM_6[31:18]};	// sequencer-master.scala:109:14
        e_0_base_vp_id = _RANDOM_8[21:18];	// sequencer-master.scala:109:14
        e_0_base_vp_valid = _RANDOM_8[22];	// sequencer-master.scala:109:14
        e_0_base_vp_scalar = _RANDOM_8[23];	// sequencer-master.scala:109:14
        e_0_base_vp_pred = _RANDOM_8[24];	// sequencer-master.scala:109:14
        _RANDOM_9 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_base_vs1_id = {_RANDOM_9[0], _RANDOM_8[31:25]};	// sequencer-master.scala:109:14
        e_0_base_vs1_valid = _RANDOM_9[1];	// sequencer-master.scala:109:14
        e_0_base_vs1_scalar = _RANDOM_9[2];	// sequencer-master.scala:109:14
        e_0_base_vs1_pred = _RANDOM_9[3];	// sequencer-master.scala:109:14
        e_0_base_vs1_prec = _RANDOM_9[5:4];	// sequencer-master.scala:109:14
        e_0_base_vs2_id = _RANDOM_9[13:6];	// sequencer-master.scala:109:14
        e_0_base_vs2_valid = _RANDOM_9[14];	// sequencer-master.scala:109:14
        e_0_base_vs2_scalar = _RANDOM_9[15];	// sequencer-master.scala:109:14
        e_0_base_vs2_pred = _RANDOM_9[16];	// sequencer-master.scala:109:14
        e_0_base_vs2_prec = _RANDOM_9[18:17];	// sequencer-master.scala:109:14
        e_0_base_vs3_id = _RANDOM_9[26:19];	// sequencer-master.scala:109:14
        e_0_base_vs3_valid = _RANDOM_9[27];	// sequencer-master.scala:109:14
        e_0_base_vs3_scalar = _RANDOM_9[28];	// sequencer-master.scala:109:14
        e_0_base_vs3_pred = _RANDOM_9[29];	// sequencer-master.scala:109:14
        e_0_base_vs3_prec = _RANDOM_9[31:30];	// sequencer-master.scala:109:14
        _RANDOM_10 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_base_vd_id = _RANDOM_10[7:0];	// sequencer-master.scala:109:14
        e_0_base_vd_valid = _RANDOM_10[8];	// sequencer-master.scala:109:14
        e_0_base_vd_scalar = _RANDOM_10[9];	// sequencer-master.scala:109:14
        e_0_base_vd_pred = _RANDOM_10[10];	// sequencer-master.scala:109:14
        e_0_base_vd_prec = _RANDOM_10[12:11];	// sequencer-master.scala:109:14
        e_0_active_viu = _RANDOM_10[13];	// sequencer-master.scala:109:14
        e_0_active_vipu = _RANDOM_10[14];	// sequencer-master.scala:109:14
        e_0_active_vimu = _RANDOM_10[15];	// sequencer-master.scala:109:14
        e_0_active_vidu = _RANDOM_10[16];	// sequencer-master.scala:109:14
        e_0_active_vfmu = _RANDOM_10[17];	// sequencer-master.scala:109:14
        e_0_active_vfdu = _RANDOM_10[18];	// sequencer-master.scala:109:14
        e_0_active_vfcu = _RANDOM_10[19];	// sequencer-master.scala:109:14
        e_0_active_vfvu = _RANDOM_10[20];	// sequencer-master.scala:109:14
        e_0_active_vpu = _RANDOM_10[21];	// sequencer-master.scala:109:14
        e_0_active_vgu = _RANDOM_10[22];	// sequencer-master.scala:109:14
        e_0_active_vcu = _RANDOM_10[23];	// sequencer-master.scala:109:14
        e_0_active_vlu = _RANDOM_10[24];	// sequencer-master.scala:109:14
        e_0_active_vsu = _RANDOM_10[25];	// sequencer-master.scala:109:14
        e_0_active_vqu = _RANDOM_10[26];	// sequencer-master.scala:109:14
        e_0_raw_0 = _RANDOM_10[27];	// sequencer-master.scala:109:14
        e_0_raw_1 = _RANDOM_10[28];	// sequencer-master.scala:109:14
        e_0_raw_2 = _RANDOM_10[29];	// sequencer-master.scala:109:14
        e_0_raw_3 = _RANDOM_10[30];	// sequencer-master.scala:109:14
        e_0_raw_4 = _RANDOM_10[31];	// sequencer-master.scala:109:14
        _RANDOM_11 = `RANDOM;	// sequencer-master.scala:109:14
        e_0_raw_5 = _RANDOM_11[0];	// sequencer-master.scala:109:14
        e_0_raw_6 = _RANDOM_11[1];	// sequencer-master.scala:109:14
        e_0_raw_7 = _RANDOM_11[2];	// sequencer-master.scala:109:14
        e_0_war_0 = _RANDOM_11[3];	// sequencer-master.scala:109:14
        e_0_war_1 = _RANDOM_11[4];	// sequencer-master.scala:109:14
        e_0_war_2 = _RANDOM_11[5];	// sequencer-master.scala:109:14
        e_0_war_3 = _RANDOM_11[6];	// sequencer-master.scala:109:14
        e_0_war_4 = _RANDOM_11[7];	// sequencer-master.scala:109:14
        e_0_war_5 = _RANDOM_11[8];	// sequencer-master.scala:109:14
        e_0_war_6 = _RANDOM_11[9];	// sequencer-master.scala:109:14
        e_0_war_7 = _RANDOM_11[10];	// sequencer-master.scala:109:14
        e_0_waw_0 = _RANDOM_11[11];	// sequencer-master.scala:109:14
        e_0_waw_1 = _RANDOM_11[12];	// sequencer-master.scala:109:14
        e_0_waw_2 = _RANDOM_11[13];	// sequencer-master.scala:109:14
        e_0_waw_3 = _RANDOM_11[14];	// sequencer-master.scala:109:14
        e_0_waw_4 = _RANDOM_11[15];	// sequencer-master.scala:109:14
        e_0_waw_5 = _RANDOM_11[16];	// sequencer-master.scala:109:14
        e_0_waw_6 = _RANDOM_11[17];	// sequencer-master.scala:109:14
        e_0_waw_7 = _RANDOM_11[18];	// sequencer-master.scala:109:14
        e_0_last = _RANDOM_11[19];	// sequencer-master.scala:109:14
        e_0_rports = _RANDOM_11[21:20];	// sequencer-master.scala:109:14
        e_0_wport_sram = _RANDOM_11[25:22];	// sequencer-master.scala:109:14
        e_0_wport_pred = _RANDOM_11[28:26];	// sequencer-master.scala:109:14
        _RANDOM_12 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_fn_union = {_RANDOM_12[6:0], _RANDOM_11[31:29]};	// sequencer-master.scala:109:14
        _RANDOM_13 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_14 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_sreg_ss1 = {_RANDOM_14[6:0], _RANDOM_13, _RANDOM_12[31:7]};	// sequencer-master.scala:109:14
        _RANDOM_15 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_16 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_sreg_ss2 = {_RANDOM_16[6:0], _RANDOM_15, _RANDOM_14[31:7]};	// sequencer-master.scala:109:14
        _RANDOM_17 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_18 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_sreg_ss3 = {_RANDOM_18[6:0], _RANDOM_17, _RANDOM_16[31:7]};	// sequencer-master.scala:109:14
        e_1_base_vp_id = _RANDOM_18[10:7];	// sequencer-master.scala:109:14
        e_1_base_vp_valid = _RANDOM_18[11];	// sequencer-master.scala:109:14
        e_1_base_vp_scalar = _RANDOM_18[12];	// sequencer-master.scala:109:14
        e_1_base_vp_pred = _RANDOM_18[13];	// sequencer-master.scala:109:14
        e_1_base_vs1_id = _RANDOM_18[21:14];	// sequencer-master.scala:109:14
        e_1_base_vs1_valid = _RANDOM_18[22];	// sequencer-master.scala:109:14
        e_1_base_vs1_scalar = _RANDOM_18[23];	// sequencer-master.scala:109:14
        e_1_base_vs1_pred = _RANDOM_18[24];	// sequencer-master.scala:109:14
        e_1_base_vs1_prec = _RANDOM_18[26:25];	// sequencer-master.scala:109:14
        _RANDOM_19 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_base_vs2_id = {_RANDOM_19[2:0], _RANDOM_18[31:27]};	// sequencer-master.scala:109:14
        e_1_base_vs2_valid = _RANDOM_19[3];	// sequencer-master.scala:109:14
        e_1_base_vs2_scalar = _RANDOM_19[4];	// sequencer-master.scala:109:14
        e_1_base_vs2_pred = _RANDOM_19[5];	// sequencer-master.scala:109:14
        e_1_base_vs2_prec = _RANDOM_19[7:6];	// sequencer-master.scala:109:14
        e_1_base_vs3_id = _RANDOM_19[15:8];	// sequencer-master.scala:109:14
        e_1_base_vs3_valid = _RANDOM_19[16];	// sequencer-master.scala:109:14
        e_1_base_vs3_scalar = _RANDOM_19[17];	// sequencer-master.scala:109:14
        e_1_base_vs3_pred = _RANDOM_19[18];	// sequencer-master.scala:109:14
        e_1_base_vs3_prec = _RANDOM_19[20:19];	// sequencer-master.scala:109:14
        e_1_base_vd_id = _RANDOM_19[28:21];	// sequencer-master.scala:109:14
        e_1_base_vd_valid = _RANDOM_19[29];	// sequencer-master.scala:109:14
        e_1_base_vd_scalar = _RANDOM_19[30];	// sequencer-master.scala:109:14
        e_1_base_vd_pred = _RANDOM_19[31];	// sequencer-master.scala:109:14
        _RANDOM_20 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_base_vd_prec = _RANDOM_20[1:0];	// sequencer-master.scala:109:14
        e_1_active_viu = _RANDOM_20[2];	// sequencer-master.scala:109:14
        e_1_active_vipu = _RANDOM_20[3];	// sequencer-master.scala:109:14
        e_1_active_vimu = _RANDOM_20[4];	// sequencer-master.scala:109:14
        e_1_active_vidu = _RANDOM_20[5];	// sequencer-master.scala:109:14
        e_1_active_vfmu = _RANDOM_20[6];	// sequencer-master.scala:109:14
        e_1_active_vfdu = _RANDOM_20[7];	// sequencer-master.scala:109:14
        e_1_active_vfcu = _RANDOM_20[8];	// sequencer-master.scala:109:14
        e_1_active_vfvu = _RANDOM_20[9];	// sequencer-master.scala:109:14
        e_1_active_vpu = _RANDOM_20[10];	// sequencer-master.scala:109:14
        e_1_active_vgu = _RANDOM_20[11];	// sequencer-master.scala:109:14
        e_1_active_vcu = _RANDOM_20[12];	// sequencer-master.scala:109:14
        e_1_active_vlu = _RANDOM_20[13];	// sequencer-master.scala:109:14
        e_1_active_vsu = _RANDOM_20[14];	// sequencer-master.scala:109:14
        e_1_active_vqu = _RANDOM_20[15];	// sequencer-master.scala:109:14
        e_1_raw_0 = _RANDOM_20[16];	// sequencer-master.scala:109:14
        e_1_raw_1 = _RANDOM_20[17];	// sequencer-master.scala:109:14
        e_1_raw_2 = _RANDOM_20[18];	// sequencer-master.scala:109:14
        e_1_raw_3 = _RANDOM_20[19];	// sequencer-master.scala:109:14
        e_1_raw_4 = _RANDOM_20[20];	// sequencer-master.scala:109:14
        e_1_raw_5 = _RANDOM_20[21];	// sequencer-master.scala:109:14
        e_1_raw_6 = _RANDOM_20[22];	// sequencer-master.scala:109:14
        e_1_raw_7 = _RANDOM_20[23];	// sequencer-master.scala:109:14
        e_1_war_0 = _RANDOM_20[24];	// sequencer-master.scala:109:14
        e_1_war_1 = _RANDOM_20[25];	// sequencer-master.scala:109:14
        e_1_war_2 = _RANDOM_20[26];	// sequencer-master.scala:109:14
        e_1_war_3 = _RANDOM_20[27];	// sequencer-master.scala:109:14
        e_1_war_4 = _RANDOM_20[28];	// sequencer-master.scala:109:14
        e_1_war_5 = _RANDOM_20[29];	// sequencer-master.scala:109:14
        e_1_war_6 = _RANDOM_20[30];	// sequencer-master.scala:109:14
        e_1_war_7 = _RANDOM_20[31];	// sequencer-master.scala:109:14
        _RANDOM_21 = `RANDOM;	// sequencer-master.scala:109:14
        e_1_waw_0 = _RANDOM_21[0];	// sequencer-master.scala:109:14
        e_1_waw_1 = _RANDOM_21[1];	// sequencer-master.scala:109:14
        e_1_waw_2 = _RANDOM_21[2];	// sequencer-master.scala:109:14
        e_1_waw_3 = _RANDOM_21[3];	// sequencer-master.scala:109:14
        e_1_waw_4 = _RANDOM_21[4];	// sequencer-master.scala:109:14
        e_1_waw_5 = _RANDOM_21[5];	// sequencer-master.scala:109:14
        e_1_waw_6 = _RANDOM_21[6];	// sequencer-master.scala:109:14
        e_1_waw_7 = _RANDOM_21[7];	// sequencer-master.scala:109:14
        e_1_last = _RANDOM_21[8];	// sequencer-master.scala:109:14
        e_1_rports = _RANDOM_21[10:9];	// sequencer-master.scala:109:14
        e_1_wport_sram = _RANDOM_21[14:11];	// sequencer-master.scala:109:14
        e_1_wport_pred = _RANDOM_21[17:15];	// sequencer-master.scala:109:14
        e_2_fn_union = _RANDOM_21[27:18];	// sequencer-master.scala:109:14
        _RANDOM_22 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_23 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_sreg_ss1 = {_RANDOM_23[27:0], _RANDOM_22, _RANDOM_21[31:28]};	// sequencer-master.scala:109:14
        _RANDOM_24 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_25 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_sreg_ss2 = {_RANDOM_25[27:0], _RANDOM_24, _RANDOM_23[31:28]};	// sequencer-master.scala:109:14
        _RANDOM_26 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_27 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_sreg_ss3 = {_RANDOM_27[27:0], _RANDOM_26, _RANDOM_25[31:28]};	// sequencer-master.scala:109:14
        e_2_base_vp_id = _RANDOM_27[31:28];	// sequencer-master.scala:109:14
        _RANDOM_28 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_base_vp_valid = _RANDOM_28[0];	// sequencer-master.scala:109:14
        e_2_base_vp_scalar = _RANDOM_28[1];	// sequencer-master.scala:109:14
        e_2_base_vp_pred = _RANDOM_28[2];	// sequencer-master.scala:109:14
        e_2_base_vs1_id = _RANDOM_28[10:3];	// sequencer-master.scala:109:14
        e_2_base_vs1_valid = _RANDOM_28[11];	// sequencer-master.scala:109:14
        e_2_base_vs1_scalar = _RANDOM_28[12];	// sequencer-master.scala:109:14
        e_2_base_vs1_pred = _RANDOM_28[13];	// sequencer-master.scala:109:14
        e_2_base_vs1_prec = _RANDOM_28[15:14];	// sequencer-master.scala:109:14
        e_2_base_vs2_id = _RANDOM_28[23:16];	// sequencer-master.scala:109:14
        e_2_base_vs2_valid = _RANDOM_28[24];	// sequencer-master.scala:109:14
        e_2_base_vs2_scalar = _RANDOM_28[25];	// sequencer-master.scala:109:14
        e_2_base_vs2_pred = _RANDOM_28[26];	// sequencer-master.scala:109:14
        e_2_base_vs2_prec = _RANDOM_28[28:27];	// sequencer-master.scala:109:14
        _RANDOM_29 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_base_vs3_id = {_RANDOM_29[4:0], _RANDOM_28[31:29]};	// sequencer-master.scala:109:14
        e_2_base_vs3_valid = _RANDOM_29[5];	// sequencer-master.scala:109:14
        e_2_base_vs3_scalar = _RANDOM_29[6];	// sequencer-master.scala:109:14
        e_2_base_vs3_pred = _RANDOM_29[7];	// sequencer-master.scala:109:14
        e_2_base_vs3_prec = _RANDOM_29[9:8];	// sequencer-master.scala:109:14
        e_2_base_vd_id = _RANDOM_29[17:10];	// sequencer-master.scala:109:14
        e_2_base_vd_valid = _RANDOM_29[18];	// sequencer-master.scala:109:14
        e_2_base_vd_scalar = _RANDOM_29[19];	// sequencer-master.scala:109:14
        e_2_base_vd_pred = _RANDOM_29[20];	// sequencer-master.scala:109:14
        e_2_base_vd_prec = _RANDOM_29[22:21];	// sequencer-master.scala:109:14
        e_2_active_viu = _RANDOM_29[23];	// sequencer-master.scala:109:14
        e_2_active_vipu = _RANDOM_29[24];	// sequencer-master.scala:109:14
        e_2_active_vimu = _RANDOM_29[25];	// sequencer-master.scala:109:14
        e_2_active_vidu = _RANDOM_29[26];	// sequencer-master.scala:109:14
        e_2_active_vfmu = _RANDOM_29[27];	// sequencer-master.scala:109:14
        e_2_active_vfdu = _RANDOM_29[28];	// sequencer-master.scala:109:14
        e_2_active_vfcu = _RANDOM_29[29];	// sequencer-master.scala:109:14
        e_2_active_vfvu = _RANDOM_29[30];	// sequencer-master.scala:109:14
        e_2_active_vpu = _RANDOM_29[31];	// sequencer-master.scala:109:14
        _RANDOM_30 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_active_vgu = _RANDOM_30[0];	// sequencer-master.scala:109:14
        e_2_active_vcu = _RANDOM_30[1];	// sequencer-master.scala:109:14
        e_2_active_vlu = _RANDOM_30[2];	// sequencer-master.scala:109:14
        e_2_active_vsu = _RANDOM_30[3];	// sequencer-master.scala:109:14
        e_2_active_vqu = _RANDOM_30[4];	// sequencer-master.scala:109:14
        e_2_raw_0 = _RANDOM_30[5];	// sequencer-master.scala:109:14
        e_2_raw_1 = _RANDOM_30[6];	// sequencer-master.scala:109:14
        e_2_raw_2 = _RANDOM_30[7];	// sequencer-master.scala:109:14
        e_2_raw_3 = _RANDOM_30[8];	// sequencer-master.scala:109:14
        e_2_raw_4 = _RANDOM_30[9];	// sequencer-master.scala:109:14
        e_2_raw_5 = _RANDOM_30[10];	// sequencer-master.scala:109:14
        e_2_raw_6 = _RANDOM_30[11];	// sequencer-master.scala:109:14
        e_2_raw_7 = _RANDOM_30[12];	// sequencer-master.scala:109:14
        e_2_war_0 = _RANDOM_30[13];	// sequencer-master.scala:109:14
        e_2_war_1 = _RANDOM_30[14];	// sequencer-master.scala:109:14
        e_2_war_2 = _RANDOM_30[15];	// sequencer-master.scala:109:14
        e_2_war_3 = _RANDOM_30[16];	// sequencer-master.scala:109:14
        e_2_war_4 = _RANDOM_30[17];	// sequencer-master.scala:109:14
        e_2_war_5 = _RANDOM_30[18];	// sequencer-master.scala:109:14
        e_2_war_6 = _RANDOM_30[19];	// sequencer-master.scala:109:14
        e_2_war_7 = _RANDOM_30[20];	// sequencer-master.scala:109:14
        e_2_waw_0 = _RANDOM_30[21];	// sequencer-master.scala:109:14
        e_2_waw_1 = _RANDOM_30[22];	// sequencer-master.scala:109:14
        e_2_waw_2 = _RANDOM_30[23];	// sequencer-master.scala:109:14
        e_2_waw_3 = _RANDOM_30[24];	// sequencer-master.scala:109:14
        e_2_waw_4 = _RANDOM_30[25];	// sequencer-master.scala:109:14
        e_2_waw_5 = _RANDOM_30[26];	// sequencer-master.scala:109:14
        e_2_waw_6 = _RANDOM_30[27];	// sequencer-master.scala:109:14
        e_2_waw_7 = _RANDOM_30[28];	// sequencer-master.scala:109:14
        e_2_last = _RANDOM_30[29];	// sequencer-master.scala:109:14
        e_2_rports = _RANDOM_30[31:30];	// sequencer-master.scala:109:14
        _RANDOM_31 = `RANDOM;	// sequencer-master.scala:109:14
        e_2_wport_sram = _RANDOM_31[3:0];	// sequencer-master.scala:109:14
        e_2_wport_pred = _RANDOM_31[6:4];	// sequencer-master.scala:109:14
        e_3_fn_union = _RANDOM_31[16:7];	// sequencer-master.scala:109:14
        _RANDOM_32 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_33 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_sreg_ss1 = {_RANDOM_33[16:0], _RANDOM_32, _RANDOM_31[31:17]};	// sequencer-master.scala:109:14
        _RANDOM_34 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_35 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_sreg_ss2 = {_RANDOM_35[16:0], _RANDOM_34, _RANDOM_33[31:17]};	// sequencer-master.scala:109:14
        _RANDOM_36 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_37 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_sreg_ss3 = {_RANDOM_37[16:0], _RANDOM_36, _RANDOM_35[31:17]};	// sequencer-master.scala:109:14
        e_3_base_vp_id = _RANDOM_37[20:17];	// sequencer-master.scala:109:14
        e_3_base_vp_valid = _RANDOM_37[21];	// sequencer-master.scala:109:14
        e_3_base_vp_scalar = _RANDOM_37[22];	// sequencer-master.scala:109:14
        e_3_base_vp_pred = _RANDOM_37[23];	// sequencer-master.scala:109:14
        e_3_base_vs1_id = _RANDOM_37[31:24];	// sequencer-master.scala:109:14
        _RANDOM_38 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_base_vs1_valid = _RANDOM_38[0];	// sequencer-master.scala:109:14
        e_3_base_vs1_scalar = _RANDOM_38[1];	// sequencer-master.scala:109:14
        e_3_base_vs1_pred = _RANDOM_38[2];	// sequencer-master.scala:109:14
        e_3_base_vs1_prec = _RANDOM_38[4:3];	// sequencer-master.scala:109:14
        e_3_base_vs2_id = _RANDOM_38[12:5];	// sequencer-master.scala:109:14
        e_3_base_vs2_valid = _RANDOM_38[13];	// sequencer-master.scala:109:14
        e_3_base_vs2_scalar = _RANDOM_38[14];	// sequencer-master.scala:109:14
        e_3_base_vs2_pred = _RANDOM_38[15];	// sequencer-master.scala:109:14
        e_3_base_vs2_prec = _RANDOM_38[17:16];	// sequencer-master.scala:109:14
        e_3_base_vs3_id = _RANDOM_38[25:18];	// sequencer-master.scala:109:14
        e_3_base_vs3_valid = _RANDOM_38[26];	// sequencer-master.scala:109:14
        e_3_base_vs3_scalar = _RANDOM_38[27];	// sequencer-master.scala:109:14
        e_3_base_vs3_pred = _RANDOM_38[28];	// sequencer-master.scala:109:14
        e_3_base_vs3_prec = _RANDOM_38[30:29];	// sequencer-master.scala:109:14
        _RANDOM_39 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_base_vd_id = {_RANDOM_39[6:0], _RANDOM_38[31]};	// sequencer-master.scala:109:14
        e_3_base_vd_valid = _RANDOM_39[7];	// sequencer-master.scala:109:14
        e_3_base_vd_scalar = _RANDOM_39[8];	// sequencer-master.scala:109:14
        e_3_base_vd_pred = _RANDOM_39[9];	// sequencer-master.scala:109:14
        e_3_base_vd_prec = _RANDOM_39[11:10];	// sequencer-master.scala:109:14
        e_3_active_viu = _RANDOM_39[12];	// sequencer-master.scala:109:14
        e_3_active_vipu = _RANDOM_39[13];	// sequencer-master.scala:109:14
        e_3_active_vimu = _RANDOM_39[14];	// sequencer-master.scala:109:14
        e_3_active_vidu = _RANDOM_39[15];	// sequencer-master.scala:109:14
        e_3_active_vfmu = _RANDOM_39[16];	// sequencer-master.scala:109:14
        e_3_active_vfdu = _RANDOM_39[17];	// sequencer-master.scala:109:14
        e_3_active_vfcu = _RANDOM_39[18];	// sequencer-master.scala:109:14
        e_3_active_vfvu = _RANDOM_39[19];	// sequencer-master.scala:109:14
        e_3_active_vpu = _RANDOM_39[20];	// sequencer-master.scala:109:14
        e_3_active_vgu = _RANDOM_39[21];	// sequencer-master.scala:109:14
        e_3_active_vcu = _RANDOM_39[22];	// sequencer-master.scala:109:14
        e_3_active_vlu = _RANDOM_39[23];	// sequencer-master.scala:109:14
        e_3_active_vsu = _RANDOM_39[24];	// sequencer-master.scala:109:14
        e_3_active_vqu = _RANDOM_39[25];	// sequencer-master.scala:109:14
        e_3_raw_0 = _RANDOM_39[26];	// sequencer-master.scala:109:14
        e_3_raw_1 = _RANDOM_39[27];	// sequencer-master.scala:109:14
        e_3_raw_2 = _RANDOM_39[28];	// sequencer-master.scala:109:14
        e_3_raw_3 = _RANDOM_39[29];	// sequencer-master.scala:109:14
        e_3_raw_4 = _RANDOM_39[30];	// sequencer-master.scala:109:14
        e_3_raw_5 = _RANDOM_39[31];	// sequencer-master.scala:109:14
        _RANDOM_40 = `RANDOM;	// sequencer-master.scala:109:14
        e_3_raw_6 = _RANDOM_40[0];	// sequencer-master.scala:109:14
        e_3_raw_7 = _RANDOM_40[1];	// sequencer-master.scala:109:14
        e_3_war_0 = _RANDOM_40[2];	// sequencer-master.scala:109:14
        e_3_war_1 = _RANDOM_40[3];	// sequencer-master.scala:109:14
        e_3_war_2 = _RANDOM_40[4];	// sequencer-master.scala:109:14
        e_3_war_3 = _RANDOM_40[5];	// sequencer-master.scala:109:14
        e_3_war_4 = _RANDOM_40[6];	// sequencer-master.scala:109:14
        e_3_war_5 = _RANDOM_40[7];	// sequencer-master.scala:109:14
        e_3_war_6 = _RANDOM_40[8];	// sequencer-master.scala:109:14
        e_3_war_7 = _RANDOM_40[9];	// sequencer-master.scala:109:14
        e_3_waw_0 = _RANDOM_40[10];	// sequencer-master.scala:109:14
        e_3_waw_1 = _RANDOM_40[11];	// sequencer-master.scala:109:14
        e_3_waw_2 = _RANDOM_40[12];	// sequencer-master.scala:109:14
        e_3_waw_3 = _RANDOM_40[13];	// sequencer-master.scala:109:14
        e_3_waw_4 = _RANDOM_40[14];	// sequencer-master.scala:109:14
        e_3_waw_5 = _RANDOM_40[15];	// sequencer-master.scala:109:14
        e_3_waw_6 = _RANDOM_40[16];	// sequencer-master.scala:109:14
        e_3_waw_7 = _RANDOM_40[17];	// sequencer-master.scala:109:14
        e_3_last = _RANDOM_40[18];	// sequencer-master.scala:109:14
        e_3_rports = _RANDOM_40[20:19];	// sequencer-master.scala:109:14
        e_3_wport_sram = _RANDOM_40[24:21];	// sequencer-master.scala:109:14
        e_3_wport_pred = _RANDOM_40[27:25];	// sequencer-master.scala:109:14
        _RANDOM_41 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_fn_union = {_RANDOM_41[5:0], _RANDOM_40[31:28]};	// sequencer-master.scala:109:14
        _RANDOM_42 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_43 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_sreg_ss1 = {_RANDOM_43[5:0], _RANDOM_42, _RANDOM_41[31:6]};	// sequencer-master.scala:109:14
        _RANDOM_44 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_45 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_sreg_ss2 = {_RANDOM_45[5:0], _RANDOM_44, _RANDOM_43[31:6]};	// sequencer-master.scala:109:14
        _RANDOM_46 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_47 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_sreg_ss3 = {_RANDOM_47[5:0], _RANDOM_46, _RANDOM_45[31:6]};	// sequencer-master.scala:109:14
        e_4_base_vp_id = _RANDOM_47[9:6];	// sequencer-master.scala:109:14
        e_4_base_vp_valid = _RANDOM_47[10];	// sequencer-master.scala:109:14
        e_4_base_vp_scalar = _RANDOM_47[11];	// sequencer-master.scala:109:14
        e_4_base_vp_pred = _RANDOM_47[12];	// sequencer-master.scala:109:14
        e_4_base_vs1_id = _RANDOM_47[20:13];	// sequencer-master.scala:109:14
        e_4_base_vs1_valid = _RANDOM_47[21];	// sequencer-master.scala:109:14
        e_4_base_vs1_scalar = _RANDOM_47[22];	// sequencer-master.scala:109:14
        e_4_base_vs1_pred = _RANDOM_47[23];	// sequencer-master.scala:109:14
        e_4_base_vs1_prec = _RANDOM_47[25:24];	// sequencer-master.scala:109:14
        _RANDOM_48 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_base_vs2_id = {_RANDOM_48[1:0], _RANDOM_47[31:26]};	// sequencer-master.scala:109:14
        e_4_base_vs2_valid = _RANDOM_48[2];	// sequencer-master.scala:109:14
        e_4_base_vs2_scalar = _RANDOM_48[3];	// sequencer-master.scala:109:14
        e_4_base_vs2_pred = _RANDOM_48[4];	// sequencer-master.scala:109:14
        e_4_base_vs2_prec = _RANDOM_48[6:5];	// sequencer-master.scala:109:14
        e_4_base_vs3_id = _RANDOM_48[14:7];	// sequencer-master.scala:109:14
        e_4_base_vs3_valid = _RANDOM_48[15];	// sequencer-master.scala:109:14
        e_4_base_vs3_scalar = _RANDOM_48[16];	// sequencer-master.scala:109:14
        e_4_base_vs3_pred = _RANDOM_48[17];	// sequencer-master.scala:109:14
        e_4_base_vs3_prec = _RANDOM_48[19:18];	// sequencer-master.scala:109:14
        e_4_base_vd_id = _RANDOM_48[27:20];	// sequencer-master.scala:109:14
        e_4_base_vd_valid = _RANDOM_48[28];	// sequencer-master.scala:109:14
        e_4_base_vd_scalar = _RANDOM_48[29];	// sequencer-master.scala:109:14
        e_4_base_vd_pred = _RANDOM_48[30];	// sequencer-master.scala:109:14
        _RANDOM_49 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_base_vd_prec = {_RANDOM_49[0], _RANDOM_48[31]};	// sequencer-master.scala:109:14
        e_4_active_viu = _RANDOM_49[1];	// sequencer-master.scala:109:14
        e_4_active_vipu = _RANDOM_49[2];	// sequencer-master.scala:109:14
        e_4_active_vimu = _RANDOM_49[3];	// sequencer-master.scala:109:14
        e_4_active_vidu = _RANDOM_49[4];	// sequencer-master.scala:109:14
        e_4_active_vfmu = _RANDOM_49[5];	// sequencer-master.scala:109:14
        e_4_active_vfdu = _RANDOM_49[6];	// sequencer-master.scala:109:14
        e_4_active_vfcu = _RANDOM_49[7];	// sequencer-master.scala:109:14
        e_4_active_vfvu = _RANDOM_49[8];	// sequencer-master.scala:109:14
        e_4_active_vpu = _RANDOM_49[9];	// sequencer-master.scala:109:14
        e_4_active_vgu = _RANDOM_49[10];	// sequencer-master.scala:109:14
        e_4_active_vcu = _RANDOM_49[11];	// sequencer-master.scala:109:14
        e_4_active_vlu = _RANDOM_49[12];	// sequencer-master.scala:109:14
        e_4_active_vsu = _RANDOM_49[13];	// sequencer-master.scala:109:14
        e_4_active_vqu = _RANDOM_49[14];	// sequencer-master.scala:109:14
        e_4_raw_0 = _RANDOM_49[15];	// sequencer-master.scala:109:14
        e_4_raw_1 = _RANDOM_49[16];	// sequencer-master.scala:109:14
        e_4_raw_2 = _RANDOM_49[17];	// sequencer-master.scala:109:14
        e_4_raw_3 = _RANDOM_49[18];	// sequencer-master.scala:109:14
        e_4_raw_4 = _RANDOM_49[19];	// sequencer-master.scala:109:14
        e_4_raw_5 = _RANDOM_49[20];	// sequencer-master.scala:109:14
        e_4_raw_6 = _RANDOM_49[21];	// sequencer-master.scala:109:14
        e_4_raw_7 = _RANDOM_49[22];	// sequencer-master.scala:109:14
        e_4_war_0 = _RANDOM_49[23];	// sequencer-master.scala:109:14
        e_4_war_1 = _RANDOM_49[24];	// sequencer-master.scala:109:14
        e_4_war_2 = _RANDOM_49[25];	// sequencer-master.scala:109:14
        e_4_war_3 = _RANDOM_49[26];	// sequencer-master.scala:109:14
        e_4_war_4 = _RANDOM_49[27];	// sequencer-master.scala:109:14
        e_4_war_5 = _RANDOM_49[28];	// sequencer-master.scala:109:14
        e_4_war_6 = _RANDOM_49[29];	// sequencer-master.scala:109:14
        e_4_war_7 = _RANDOM_49[30];	// sequencer-master.scala:109:14
        e_4_waw_0 = _RANDOM_49[31];	// sequencer-master.scala:109:14
        _RANDOM_50 = `RANDOM;	// sequencer-master.scala:109:14
        e_4_waw_1 = _RANDOM_50[0];	// sequencer-master.scala:109:14
        e_4_waw_2 = _RANDOM_50[1];	// sequencer-master.scala:109:14
        e_4_waw_3 = _RANDOM_50[2];	// sequencer-master.scala:109:14
        e_4_waw_4 = _RANDOM_50[3];	// sequencer-master.scala:109:14
        e_4_waw_5 = _RANDOM_50[4];	// sequencer-master.scala:109:14
        e_4_waw_6 = _RANDOM_50[5];	// sequencer-master.scala:109:14
        e_4_waw_7 = _RANDOM_50[6];	// sequencer-master.scala:109:14
        e_4_last = _RANDOM_50[7];	// sequencer-master.scala:109:14
        e_4_rports = _RANDOM_50[9:8];	// sequencer-master.scala:109:14
        e_4_wport_sram = _RANDOM_50[13:10];	// sequencer-master.scala:109:14
        e_4_wport_pred = _RANDOM_50[16:14];	// sequencer-master.scala:109:14
        e_5_fn_union = _RANDOM_50[26:17];	// sequencer-master.scala:109:14
        _RANDOM_51 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_52 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_sreg_ss1 = {_RANDOM_52[26:0], _RANDOM_51, _RANDOM_50[31:27]};	// sequencer-master.scala:109:14
        _RANDOM_53 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_54 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_sreg_ss2 = {_RANDOM_54[26:0], _RANDOM_53, _RANDOM_52[31:27]};	// sequencer-master.scala:109:14
        _RANDOM_55 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_56 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_sreg_ss3 = {_RANDOM_56[26:0], _RANDOM_55, _RANDOM_54[31:27]};	// sequencer-master.scala:109:14
        e_5_base_vp_id = _RANDOM_56[30:27];	// sequencer-master.scala:109:14
        e_5_base_vp_valid = _RANDOM_56[31];	// sequencer-master.scala:109:14
        _RANDOM_57 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_base_vp_scalar = _RANDOM_57[0];	// sequencer-master.scala:109:14
        e_5_base_vp_pred = _RANDOM_57[1];	// sequencer-master.scala:109:14
        e_5_base_vs1_id = _RANDOM_57[9:2];	// sequencer-master.scala:109:14
        e_5_base_vs1_valid = _RANDOM_57[10];	// sequencer-master.scala:109:14
        e_5_base_vs1_scalar = _RANDOM_57[11];	// sequencer-master.scala:109:14
        e_5_base_vs1_pred = _RANDOM_57[12];	// sequencer-master.scala:109:14
        e_5_base_vs1_prec = _RANDOM_57[14:13];	// sequencer-master.scala:109:14
        e_5_base_vs2_id = _RANDOM_57[22:15];	// sequencer-master.scala:109:14
        e_5_base_vs2_valid = _RANDOM_57[23];	// sequencer-master.scala:109:14
        e_5_base_vs2_scalar = _RANDOM_57[24];	// sequencer-master.scala:109:14
        e_5_base_vs2_pred = _RANDOM_57[25];	// sequencer-master.scala:109:14
        e_5_base_vs2_prec = _RANDOM_57[27:26];	// sequencer-master.scala:109:14
        _RANDOM_58 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_base_vs3_id = {_RANDOM_58[3:0], _RANDOM_57[31:28]};	// sequencer-master.scala:109:14
        e_5_base_vs3_valid = _RANDOM_58[4];	// sequencer-master.scala:109:14
        e_5_base_vs3_scalar = _RANDOM_58[5];	// sequencer-master.scala:109:14
        e_5_base_vs3_pred = _RANDOM_58[6];	// sequencer-master.scala:109:14
        e_5_base_vs3_prec = _RANDOM_58[8:7];	// sequencer-master.scala:109:14
        e_5_base_vd_id = _RANDOM_58[16:9];	// sequencer-master.scala:109:14
        e_5_base_vd_valid = _RANDOM_58[17];	// sequencer-master.scala:109:14
        e_5_base_vd_scalar = _RANDOM_58[18];	// sequencer-master.scala:109:14
        e_5_base_vd_pred = _RANDOM_58[19];	// sequencer-master.scala:109:14
        e_5_base_vd_prec = _RANDOM_58[21:20];	// sequencer-master.scala:109:14
        e_5_active_viu = _RANDOM_58[22];	// sequencer-master.scala:109:14
        e_5_active_vipu = _RANDOM_58[23];	// sequencer-master.scala:109:14
        e_5_active_vimu = _RANDOM_58[24];	// sequencer-master.scala:109:14
        e_5_active_vidu = _RANDOM_58[25];	// sequencer-master.scala:109:14
        e_5_active_vfmu = _RANDOM_58[26];	// sequencer-master.scala:109:14
        e_5_active_vfdu = _RANDOM_58[27];	// sequencer-master.scala:109:14
        e_5_active_vfcu = _RANDOM_58[28];	// sequencer-master.scala:109:14
        e_5_active_vfvu = _RANDOM_58[29];	// sequencer-master.scala:109:14
        e_5_active_vpu = _RANDOM_58[30];	// sequencer-master.scala:109:14
        e_5_active_vgu = _RANDOM_58[31];	// sequencer-master.scala:109:14
        _RANDOM_59 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_active_vcu = _RANDOM_59[0];	// sequencer-master.scala:109:14
        e_5_active_vlu = _RANDOM_59[1];	// sequencer-master.scala:109:14
        e_5_active_vsu = _RANDOM_59[2];	// sequencer-master.scala:109:14
        e_5_active_vqu = _RANDOM_59[3];	// sequencer-master.scala:109:14
        e_5_raw_0 = _RANDOM_59[4];	// sequencer-master.scala:109:14
        e_5_raw_1 = _RANDOM_59[5];	// sequencer-master.scala:109:14
        e_5_raw_2 = _RANDOM_59[6];	// sequencer-master.scala:109:14
        e_5_raw_3 = _RANDOM_59[7];	// sequencer-master.scala:109:14
        e_5_raw_4 = _RANDOM_59[8];	// sequencer-master.scala:109:14
        e_5_raw_5 = _RANDOM_59[9];	// sequencer-master.scala:109:14
        e_5_raw_6 = _RANDOM_59[10];	// sequencer-master.scala:109:14
        e_5_raw_7 = _RANDOM_59[11];	// sequencer-master.scala:109:14
        e_5_war_0 = _RANDOM_59[12];	// sequencer-master.scala:109:14
        e_5_war_1 = _RANDOM_59[13];	// sequencer-master.scala:109:14
        e_5_war_2 = _RANDOM_59[14];	// sequencer-master.scala:109:14
        e_5_war_3 = _RANDOM_59[15];	// sequencer-master.scala:109:14
        e_5_war_4 = _RANDOM_59[16];	// sequencer-master.scala:109:14
        e_5_war_5 = _RANDOM_59[17];	// sequencer-master.scala:109:14
        e_5_war_6 = _RANDOM_59[18];	// sequencer-master.scala:109:14
        e_5_war_7 = _RANDOM_59[19];	// sequencer-master.scala:109:14
        e_5_waw_0 = _RANDOM_59[20];	// sequencer-master.scala:109:14
        e_5_waw_1 = _RANDOM_59[21];	// sequencer-master.scala:109:14
        e_5_waw_2 = _RANDOM_59[22];	// sequencer-master.scala:109:14
        e_5_waw_3 = _RANDOM_59[23];	// sequencer-master.scala:109:14
        e_5_waw_4 = _RANDOM_59[24];	// sequencer-master.scala:109:14
        e_5_waw_5 = _RANDOM_59[25];	// sequencer-master.scala:109:14
        e_5_waw_6 = _RANDOM_59[26];	// sequencer-master.scala:109:14
        e_5_waw_7 = _RANDOM_59[27];	// sequencer-master.scala:109:14
        e_5_last = _RANDOM_59[28];	// sequencer-master.scala:109:14
        e_5_rports = _RANDOM_59[30:29];	// sequencer-master.scala:109:14
        _RANDOM_60 = `RANDOM;	// sequencer-master.scala:109:14
        e_5_wport_sram = {_RANDOM_60[2:0], _RANDOM_59[31]};	// sequencer-master.scala:109:14
        e_5_wport_pred = _RANDOM_60[5:3];	// sequencer-master.scala:109:14
        e_6_fn_union = _RANDOM_60[15:6];	// sequencer-master.scala:109:14
        _RANDOM_61 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_62 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_sreg_ss1 = {_RANDOM_62[15:0], _RANDOM_61, _RANDOM_60[31:16]};	// sequencer-master.scala:109:14
        _RANDOM_63 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_64 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_sreg_ss2 = {_RANDOM_64[15:0], _RANDOM_63, _RANDOM_62[31:16]};	// sequencer-master.scala:109:14
        _RANDOM_65 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_66 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_sreg_ss3 = {_RANDOM_66[15:0], _RANDOM_65, _RANDOM_64[31:16]};	// sequencer-master.scala:109:14
        e_6_base_vp_id = _RANDOM_66[19:16];	// sequencer-master.scala:109:14
        e_6_base_vp_valid = _RANDOM_66[20];	// sequencer-master.scala:109:14
        e_6_base_vp_scalar = _RANDOM_66[21];	// sequencer-master.scala:109:14
        e_6_base_vp_pred = _RANDOM_66[22];	// sequencer-master.scala:109:14
        e_6_base_vs1_id = _RANDOM_66[30:23];	// sequencer-master.scala:109:14
        e_6_base_vs1_valid = _RANDOM_66[31];	// sequencer-master.scala:109:14
        _RANDOM_67 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_base_vs1_scalar = _RANDOM_67[0];	// sequencer-master.scala:109:14
        e_6_base_vs1_pred = _RANDOM_67[1];	// sequencer-master.scala:109:14
        e_6_base_vs1_prec = _RANDOM_67[3:2];	// sequencer-master.scala:109:14
        e_6_base_vs2_id = _RANDOM_67[11:4];	// sequencer-master.scala:109:14
        e_6_base_vs2_valid = _RANDOM_67[12];	// sequencer-master.scala:109:14
        e_6_base_vs2_scalar = _RANDOM_67[13];	// sequencer-master.scala:109:14
        e_6_base_vs2_pred = _RANDOM_67[14];	// sequencer-master.scala:109:14
        e_6_base_vs2_prec = _RANDOM_67[16:15];	// sequencer-master.scala:109:14
        e_6_base_vs3_id = _RANDOM_67[24:17];	// sequencer-master.scala:109:14
        e_6_base_vs3_valid = _RANDOM_67[25];	// sequencer-master.scala:109:14
        e_6_base_vs3_scalar = _RANDOM_67[26];	// sequencer-master.scala:109:14
        e_6_base_vs3_pred = _RANDOM_67[27];	// sequencer-master.scala:109:14
        e_6_base_vs3_prec = _RANDOM_67[29:28];	// sequencer-master.scala:109:14
        _RANDOM_68 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_base_vd_id = {_RANDOM_68[5:0], _RANDOM_67[31:30]};	// sequencer-master.scala:109:14
        e_6_base_vd_valid = _RANDOM_68[6];	// sequencer-master.scala:109:14
        e_6_base_vd_scalar = _RANDOM_68[7];	// sequencer-master.scala:109:14
        e_6_base_vd_pred = _RANDOM_68[8];	// sequencer-master.scala:109:14
        e_6_base_vd_prec = _RANDOM_68[10:9];	// sequencer-master.scala:109:14
        e_6_active_viu = _RANDOM_68[11];	// sequencer-master.scala:109:14
        e_6_active_vipu = _RANDOM_68[12];	// sequencer-master.scala:109:14
        e_6_active_vimu = _RANDOM_68[13];	// sequencer-master.scala:109:14
        e_6_active_vidu = _RANDOM_68[14];	// sequencer-master.scala:109:14
        e_6_active_vfmu = _RANDOM_68[15];	// sequencer-master.scala:109:14
        e_6_active_vfdu = _RANDOM_68[16];	// sequencer-master.scala:109:14
        e_6_active_vfcu = _RANDOM_68[17];	// sequencer-master.scala:109:14
        e_6_active_vfvu = _RANDOM_68[18];	// sequencer-master.scala:109:14
        e_6_active_vpu = _RANDOM_68[19];	// sequencer-master.scala:109:14
        e_6_active_vgu = _RANDOM_68[20];	// sequencer-master.scala:109:14
        e_6_active_vcu = _RANDOM_68[21];	// sequencer-master.scala:109:14
        e_6_active_vlu = _RANDOM_68[22];	// sequencer-master.scala:109:14
        e_6_active_vsu = _RANDOM_68[23];	// sequencer-master.scala:109:14
        e_6_active_vqu = _RANDOM_68[24];	// sequencer-master.scala:109:14
        e_6_raw_0 = _RANDOM_68[25];	// sequencer-master.scala:109:14
        e_6_raw_1 = _RANDOM_68[26];	// sequencer-master.scala:109:14
        e_6_raw_2 = _RANDOM_68[27];	// sequencer-master.scala:109:14
        e_6_raw_3 = _RANDOM_68[28];	// sequencer-master.scala:109:14
        e_6_raw_4 = _RANDOM_68[29];	// sequencer-master.scala:109:14
        e_6_raw_5 = _RANDOM_68[30];	// sequencer-master.scala:109:14
        e_6_raw_6 = _RANDOM_68[31];	// sequencer-master.scala:109:14
        _RANDOM_69 = `RANDOM;	// sequencer-master.scala:109:14
        e_6_raw_7 = _RANDOM_69[0];	// sequencer-master.scala:109:14
        e_6_war_0 = _RANDOM_69[1];	// sequencer-master.scala:109:14
        e_6_war_1 = _RANDOM_69[2];	// sequencer-master.scala:109:14
        e_6_war_2 = _RANDOM_69[3];	// sequencer-master.scala:109:14
        e_6_war_3 = _RANDOM_69[4];	// sequencer-master.scala:109:14
        e_6_war_4 = _RANDOM_69[5];	// sequencer-master.scala:109:14
        e_6_war_5 = _RANDOM_69[6];	// sequencer-master.scala:109:14
        e_6_war_6 = _RANDOM_69[7];	// sequencer-master.scala:109:14
        e_6_war_7 = _RANDOM_69[8];	// sequencer-master.scala:109:14
        e_6_waw_0 = _RANDOM_69[9];	// sequencer-master.scala:109:14
        e_6_waw_1 = _RANDOM_69[10];	// sequencer-master.scala:109:14
        e_6_waw_2 = _RANDOM_69[11];	// sequencer-master.scala:109:14
        e_6_waw_3 = _RANDOM_69[12];	// sequencer-master.scala:109:14
        e_6_waw_4 = _RANDOM_69[13];	// sequencer-master.scala:109:14
        e_6_waw_5 = _RANDOM_69[14];	// sequencer-master.scala:109:14
        e_6_waw_6 = _RANDOM_69[15];	// sequencer-master.scala:109:14
        e_6_waw_7 = _RANDOM_69[16];	// sequencer-master.scala:109:14
        e_6_last = _RANDOM_69[17];	// sequencer-master.scala:109:14
        e_6_rports = _RANDOM_69[19:18];	// sequencer-master.scala:109:14
        e_6_wport_sram = _RANDOM_69[23:20];	// sequencer-master.scala:109:14
        e_6_wport_pred = _RANDOM_69[26:24];	// sequencer-master.scala:109:14
        _RANDOM_70 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_fn_union = {_RANDOM_70[4:0], _RANDOM_69[31:27]};	// sequencer-master.scala:109:14
        _RANDOM_71 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_72 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_sreg_ss1 = {_RANDOM_72[4:0], _RANDOM_71, _RANDOM_70[31:5]};	// sequencer-master.scala:109:14
        _RANDOM_73 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_74 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_sreg_ss2 = {_RANDOM_74[4:0], _RANDOM_73, _RANDOM_72[31:5]};	// sequencer-master.scala:109:14
        _RANDOM_75 = `RANDOM;	// sequencer-master.scala:109:14
        _RANDOM_76 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_sreg_ss3 = {_RANDOM_76[4:0], _RANDOM_75, _RANDOM_74[31:5]};	// sequencer-master.scala:109:14
        e_7_base_vp_id = _RANDOM_76[8:5];	// sequencer-master.scala:109:14
        e_7_base_vp_valid = _RANDOM_76[9];	// sequencer-master.scala:109:14
        e_7_base_vp_scalar = _RANDOM_76[10];	// sequencer-master.scala:109:14
        e_7_base_vp_pred = _RANDOM_76[11];	// sequencer-master.scala:109:14
        e_7_base_vs1_id = _RANDOM_76[19:12];	// sequencer-master.scala:109:14
        e_7_base_vs1_valid = _RANDOM_76[20];	// sequencer-master.scala:109:14
        e_7_base_vs1_scalar = _RANDOM_76[21];	// sequencer-master.scala:109:14
        e_7_base_vs1_pred = _RANDOM_76[22];	// sequencer-master.scala:109:14
        e_7_base_vs1_prec = _RANDOM_76[24:23];	// sequencer-master.scala:109:14
        _RANDOM_77 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_base_vs2_id = {_RANDOM_77[0], _RANDOM_76[31:25]};	// sequencer-master.scala:109:14
        e_7_base_vs2_valid = _RANDOM_77[1];	// sequencer-master.scala:109:14
        e_7_base_vs2_scalar = _RANDOM_77[2];	// sequencer-master.scala:109:14
        e_7_base_vs2_pred = _RANDOM_77[3];	// sequencer-master.scala:109:14
        e_7_base_vs2_prec = _RANDOM_77[5:4];	// sequencer-master.scala:109:14
        e_7_base_vs3_id = _RANDOM_77[13:6];	// sequencer-master.scala:109:14
        e_7_base_vs3_valid = _RANDOM_77[14];	// sequencer-master.scala:109:14
        e_7_base_vs3_scalar = _RANDOM_77[15];	// sequencer-master.scala:109:14
        e_7_base_vs3_pred = _RANDOM_77[16];	// sequencer-master.scala:109:14
        e_7_base_vs3_prec = _RANDOM_77[18:17];	// sequencer-master.scala:109:14
        e_7_base_vd_id = _RANDOM_77[26:19];	// sequencer-master.scala:109:14
        e_7_base_vd_valid = _RANDOM_77[27];	// sequencer-master.scala:109:14
        e_7_base_vd_scalar = _RANDOM_77[28];	// sequencer-master.scala:109:14
        e_7_base_vd_pred = _RANDOM_77[29];	// sequencer-master.scala:109:14
        e_7_base_vd_prec = _RANDOM_77[31:30];	// sequencer-master.scala:109:14
        _RANDOM_78 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_active_viu = _RANDOM_78[0];	// sequencer-master.scala:109:14
        e_7_active_vipu = _RANDOM_78[1];	// sequencer-master.scala:109:14
        e_7_active_vimu = _RANDOM_78[2];	// sequencer-master.scala:109:14
        e_7_active_vidu = _RANDOM_78[3];	// sequencer-master.scala:109:14
        e_7_active_vfmu = _RANDOM_78[4];	// sequencer-master.scala:109:14
        e_7_active_vfdu = _RANDOM_78[5];	// sequencer-master.scala:109:14
        e_7_active_vfcu = _RANDOM_78[6];	// sequencer-master.scala:109:14
        e_7_active_vfvu = _RANDOM_78[7];	// sequencer-master.scala:109:14
        e_7_active_vpu = _RANDOM_78[8];	// sequencer-master.scala:109:14
        e_7_active_vgu = _RANDOM_78[9];	// sequencer-master.scala:109:14
        e_7_active_vcu = _RANDOM_78[10];	// sequencer-master.scala:109:14
        e_7_active_vlu = _RANDOM_78[11];	// sequencer-master.scala:109:14
        e_7_active_vsu = _RANDOM_78[12];	// sequencer-master.scala:109:14
        e_7_active_vqu = _RANDOM_78[13];	// sequencer-master.scala:109:14
        e_7_raw_0 = _RANDOM_78[14];	// sequencer-master.scala:109:14
        e_7_raw_1 = _RANDOM_78[15];	// sequencer-master.scala:109:14
        e_7_raw_2 = _RANDOM_78[16];	// sequencer-master.scala:109:14
        e_7_raw_3 = _RANDOM_78[17];	// sequencer-master.scala:109:14
        e_7_raw_4 = _RANDOM_78[18];	// sequencer-master.scala:109:14
        e_7_raw_5 = _RANDOM_78[19];	// sequencer-master.scala:109:14
        e_7_raw_6 = _RANDOM_78[20];	// sequencer-master.scala:109:14
        e_7_raw_7 = _RANDOM_78[21];	// sequencer-master.scala:109:14
        e_7_war_0 = _RANDOM_78[22];	// sequencer-master.scala:109:14
        e_7_war_1 = _RANDOM_78[23];	// sequencer-master.scala:109:14
        e_7_war_2 = _RANDOM_78[24];	// sequencer-master.scala:109:14
        e_7_war_3 = _RANDOM_78[25];	// sequencer-master.scala:109:14
        e_7_war_4 = _RANDOM_78[26];	// sequencer-master.scala:109:14
        e_7_war_5 = _RANDOM_78[27];	// sequencer-master.scala:109:14
        e_7_war_6 = _RANDOM_78[28];	// sequencer-master.scala:109:14
        e_7_war_7 = _RANDOM_78[29];	// sequencer-master.scala:109:14
        e_7_waw_0 = _RANDOM_78[30];	// sequencer-master.scala:109:14
        e_7_waw_1 = _RANDOM_78[31];	// sequencer-master.scala:109:14
        _RANDOM_79 = `RANDOM;	// sequencer-master.scala:109:14
        e_7_waw_2 = _RANDOM_79[0];	// sequencer-master.scala:109:14
        e_7_waw_3 = _RANDOM_79[1];	// sequencer-master.scala:109:14
        e_7_waw_4 = _RANDOM_79[2];	// sequencer-master.scala:109:14
        e_7_waw_5 = _RANDOM_79[3];	// sequencer-master.scala:109:14
        e_7_waw_6 = _RANDOM_79[4];	// sequencer-master.scala:109:14
        e_7_waw_7 = _RANDOM_79[5];	// sequencer-master.scala:109:14
        e_7_last = _RANDOM_79[6];	// sequencer-master.scala:109:14
        e_7_rports = _RANDOM_79[8:7];	// sequencer-master.scala:109:14
        e_7_wport_sram = _RANDOM_79[12:9];	// sequencer-master.scala:109:14
        e_7_wport_pred = _RANDOM_79[15:13];	// sequencer-master.scala:109:14
        maybe_full = _RANDOM_79[16];	// sequencer-master.scala:111:23
        head = _RANDOM_79[19:17];	// sequencer-master.scala:112:17
        tail = _RANDOM_79[22:20];	// sequencer-master.scala:113:17
        _T_2 = _RANDOM_79[23];	// sequencer-master.scala:444:24
      `endif
    end // initial
  `endif
      wire _T_399 = v_0 | v_1 | v_2 | v_3 | v_4 | v_5 | v_6 | v_7;	// sequencer-master.scala:136:44, :448:36
      wire _T_400 = _T_3 & io_op_bits_active_vidiv;	// sequencer-master.scala:643:40
      wire _T_401 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_402 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_403 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_404 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_405 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_406 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_407 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_408 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_409 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_410 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_411 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_412 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_413 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_414 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_415 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_416 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_417 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_418 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_419 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_420 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_421 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_422 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_423 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_424 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_425 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_426 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_427 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_428 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_429 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_430 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_431 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_432 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_433 = _T_3 & io_op_bits_active_vfdiv;	// sequencer-master.scala:645:40
      wire _T_434 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_435 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_436 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_437 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_438 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_439 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_440 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_441 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_442 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_443 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_444 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_445 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_446 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_447 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_448 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_449 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_450 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_451 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_452 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_453 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_454 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_455 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_456 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_457 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_458 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_459 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_460 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_461 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_462 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_463 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_464 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_465 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [7:0] _T_466 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_4 | _T_434 ?
                io_op_bits_base_vs2_id : e_0_base_vs2_id) : _T_434 ? io_op_bits_base_vs2_id :
                e_0_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_467 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_4 | _T_435 ?
                io_op_bits_base_vs2_scalar : e_0_base_vs2_scalar) : _T_435 ? io_op_bits_base_vs2_scalar :
                e_0_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_468 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_4 | _T_436 ?
                io_op_bits_base_vs2_pred : e_0_base_vs2_pred) : _T_436 ? io_op_bits_base_vs2_pred :
                e_0_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_469 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_4 | _T_437 ?
                io_op_bits_base_vs2_prec : e_0_base_vs2_prec) : _T_437 ? io_op_bits_base_vs2_prec :
                e_0_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_470 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_5 | _T_438 ?
                io_op_bits_base_vs2_id : e_1_base_vs2_id) : _T_438 ? io_op_bits_base_vs2_id :
                e_1_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_471 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_5 | _T_439 ?
                io_op_bits_base_vs2_scalar : e_1_base_vs2_scalar) : _T_439 ? io_op_bits_base_vs2_scalar :
                e_1_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_472 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_5 | _T_440 ?
                io_op_bits_base_vs2_pred : e_1_base_vs2_pred) : _T_440 ? io_op_bits_base_vs2_pred :
                e_1_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_473 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_5 | _T_441 ?
                io_op_bits_base_vs2_prec : e_1_base_vs2_prec) : _T_441 ? io_op_bits_base_vs2_prec :
                e_1_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_474 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_6 | _T_442 ?
                io_op_bits_base_vs2_id : e_2_base_vs2_id) : _T_442 ? io_op_bits_base_vs2_id :
                e_2_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_475 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_6 | _T_443 ?
                io_op_bits_base_vs2_scalar : e_2_base_vs2_scalar) : _T_443 ? io_op_bits_base_vs2_scalar :
                e_2_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_476 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_6 | _T_444 ?
                io_op_bits_base_vs2_pred : e_2_base_vs2_pred) : _T_444 ? io_op_bits_base_vs2_pred :
                e_2_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_477 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_6 | _T_445 ?
                io_op_bits_base_vs2_prec : e_2_base_vs2_prec) : _T_445 ? io_op_bits_base_vs2_prec :
                e_2_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_478 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_7 | _T_446 ?
                io_op_bits_base_vs2_id : e_3_base_vs2_id) : _T_446 ? io_op_bits_base_vs2_id :
                e_3_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_479 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_7 | _T_447 ?
                io_op_bits_base_vs2_scalar : e_3_base_vs2_scalar) : _T_447 ? io_op_bits_base_vs2_scalar :
                e_3_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_480 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_7 | _T_448 ?
                io_op_bits_base_vs2_pred : e_3_base_vs2_pred) : _T_448 ? io_op_bits_base_vs2_pred :
                e_3_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_481 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_7 | _T_449 ?
                io_op_bits_base_vs2_prec : e_3_base_vs2_prec) : _T_449 ? io_op_bits_base_vs2_prec :
                e_3_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_482 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_8 | _T_450 ?
                io_op_bits_base_vs2_id : e_4_base_vs2_id) : _T_450 ? io_op_bits_base_vs2_id :
                e_4_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_483 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_8 | _T_451 ?
                io_op_bits_base_vs2_scalar : e_4_base_vs2_scalar) : _T_451 ? io_op_bits_base_vs2_scalar :
                e_4_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_484 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_8 | _T_452 ?
                io_op_bits_base_vs2_pred : e_4_base_vs2_pred) : _T_452 ? io_op_bits_base_vs2_pred :
                e_4_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_485 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_8 | _T_453 ?
                io_op_bits_base_vs2_prec : e_4_base_vs2_prec) : _T_453 ? io_op_bits_base_vs2_prec :
                e_4_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_486 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_9 | _T_454 ?
                io_op_bits_base_vs2_id : e_5_base_vs2_id) : _T_454 ? io_op_bits_base_vs2_id :
                e_5_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_487 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_9 | _T_455 ?
                io_op_bits_base_vs2_scalar : e_5_base_vs2_scalar) : _T_455 ? io_op_bits_base_vs2_scalar :
                e_5_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_488 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_9 | _T_456 ?
                io_op_bits_base_vs2_pred : e_5_base_vs2_pred) : _T_456 ? io_op_bits_base_vs2_pred :
                e_5_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_489 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_9 | _T_457 ?
                io_op_bits_base_vs2_prec : e_5_base_vs2_prec) : _T_457 ? io_op_bits_base_vs2_prec :
                e_5_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_490 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_10 | _T_458 ?
                io_op_bits_base_vs2_id : e_6_base_vs2_id) : _T_458 ? io_op_bits_base_vs2_id :
                e_6_base_vs2_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_491 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_10 | _T_459 ?
                io_op_bits_base_vs2_scalar : e_6_base_vs2_scalar) : _T_459 ? io_op_bits_base_vs2_scalar :
                e_6_base_vs2_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_492 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_10 | _T_460 ?
                io_op_bits_base_vs2_pred : e_6_base_vs2_pred) : _T_460 ? io_op_bits_base_vs2_pred :
                e_6_base_vs2_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_493 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (_T_10 | _T_461 ?
                io_op_bits_base_vs2_prec : e_6_base_vs2_prec) : _T_461 ? io_op_bits_base_vs2_prec :
                e_6_base_vs2_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_494 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (&tail | _T_462 ?
                io_op_bits_base_vs2_id : e_7_base_vs2_id) : _T_462 ? io_op_bits_base_vs2_id :
                e_7_base_vs2_id;	// sequencer-master.scala:141:29, :267:35, :329:29, util.scala:94:11
      wire _T_495 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (&tail | _T_463 ?
                io_op_bits_base_vs2_scalar : e_7_base_vs2_scalar) : _T_463 ? io_op_bits_base_vs2_scalar :
                e_7_base_vs2_scalar;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:37, util.scala:94:11
      wire _T_496 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (&tail | _T_464 ?
                io_op_bits_base_vs2_pred : e_7_base_vs2_pred) : _T_464 ? io_op_bits_base_vs2_pred :
                e_7_base_vs2_pred;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:31, util.scala:94:11
      wire [1:0] _T_497 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid ? (&tail | _T_465 ?
                io_op_bits_base_vs2_prec : e_7_base_vs2_prec) : _T_465 ? io_op_bits_base_vs2_prec :
                e_7_base_vs2_prec;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_498 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_499 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_500 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_501 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_502 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_503 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_504 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_505 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_506 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_507 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_508 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_509 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_510 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_511 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_512 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_513 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_514 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_515 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_516 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_517 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_518 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_519 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_520 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_521 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_522 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_523 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_524 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_525 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_526 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_527 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_528 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_529 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [7:0] _T_530 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_498 ?
                io_op_bits_base_vs2_id : _T_466) : _T_498 ? io_op_bits_base_vs2_id : _T_466;	// sequencer-master.scala:329:29
      wire _T_531 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_499 ?
                io_op_bits_base_vs2_scalar : _T_467) : _T_499 ? io_op_bits_base_vs2_scalar : _T_467;	// sequencer-master.scala:329:29
      wire _T_532 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_500 ?
                io_op_bits_base_vs2_pred : _T_468) : _T_500 ? io_op_bits_base_vs2_pred : _T_468;	// sequencer-master.scala:329:29
      wire [1:0] _T_533 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_501 ?
                io_op_bits_base_vs2_prec : _T_469) : _T_501 ? io_op_bits_base_vs2_prec : _T_469;	// sequencer-master.scala:329:29
      wire [7:0] _T_534 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_502 ?
                io_op_bits_base_vs2_id : _T_470) : _T_502 ? io_op_bits_base_vs2_id : _T_470;	// sequencer-master.scala:329:29
      wire _T_535 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_503 ?
                io_op_bits_base_vs2_scalar : _T_471) : _T_503 ? io_op_bits_base_vs2_scalar : _T_471;	// sequencer-master.scala:329:29
      wire _T_536 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_504 ?
                io_op_bits_base_vs2_pred : _T_472) : _T_504 ? io_op_bits_base_vs2_pred : _T_472;	// sequencer-master.scala:329:29
      wire [1:0] _T_537 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_505 ?
                io_op_bits_base_vs2_prec : _T_473) : _T_505 ? io_op_bits_base_vs2_prec : _T_473;	// sequencer-master.scala:329:29
      wire [7:0] _T_538 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_506 ?
                io_op_bits_base_vs2_id : _T_474) : _T_506 ? io_op_bits_base_vs2_id : _T_474;	// sequencer-master.scala:329:29
      wire _T_539 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_507 ?
                io_op_bits_base_vs2_scalar : _T_475) : _T_507 ? io_op_bits_base_vs2_scalar : _T_475;	// sequencer-master.scala:329:29
      wire _T_540 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_508 ?
                io_op_bits_base_vs2_pred : _T_476) : _T_508 ? io_op_bits_base_vs2_pred : _T_476;	// sequencer-master.scala:329:29
      wire [1:0] _T_541 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_509 ?
                io_op_bits_base_vs2_prec : _T_477) : _T_509 ? io_op_bits_base_vs2_prec : _T_477;	// sequencer-master.scala:329:29
      wire [7:0] _T_542 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_510 ?
                io_op_bits_base_vs2_id : _T_478) : _T_510 ? io_op_bits_base_vs2_id : _T_478;	// sequencer-master.scala:329:29
      wire _T_543 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_511 ?
                io_op_bits_base_vs2_scalar : _T_479) : _T_511 ? io_op_bits_base_vs2_scalar : _T_479;	// sequencer-master.scala:329:29
      wire _T_544 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_512 ?
                io_op_bits_base_vs2_pred : _T_480) : _T_512 ? io_op_bits_base_vs2_pred : _T_480;	// sequencer-master.scala:329:29
      wire [1:0] _T_545 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_513 ?
                io_op_bits_base_vs2_prec : _T_481) : _T_513 ? io_op_bits_base_vs2_prec : _T_481;	// sequencer-master.scala:329:29
      wire [7:0] _T_546 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_514 ?
                io_op_bits_base_vs2_id : _T_482) : _T_514 ? io_op_bits_base_vs2_id : _T_482;	// sequencer-master.scala:329:29
      wire _T_547 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_515 ?
                io_op_bits_base_vs2_scalar : _T_483) : _T_515 ? io_op_bits_base_vs2_scalar : _T_483;	// sequencer-master.scala:329:29
      wire _T_548 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_516 ?
                io_op_bits_base_vs2_pred : _T_484) : _T_516 ? io_op_bits_base_vs2_pred : _T_484;	// sequencer-master.scala:329:29
      wire [1:0] _T_549 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_517 ?
                io_op_bits_base_vs2_prec : _T_485) : _T_517 ? io_op_bits_base_vs2_prec : _T_485;	// sequencer-master.scala:329:29
      wire [7:0] _T_550 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_518 ?
                io_op_bits_base_vs2_id : _T_486) : _T_518 ? io_op_bits_base_vs2_id : _T_486;	// sequencer-master.scala:329:29
      wire _T_551 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_519 ?
                io_op_bits_base_vs2_scalar : _T_487) : _T_519 ? io_op_bits_base_vs2_scalar : _T_487;	// sequencer-master.scala:329:29
      wire _T_552 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_520 ?
                io_op_bits_base_vs2_pred : _T_488) : _T_520 ? io_op_bits_base_vs2_pred : _T_488;	// sequencer-master.scala:329:29
      wire [1:0] _T_553 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_521 ?
                io_op_bits_base_vs2_prec : _T_489) : _T_521 ? io_op_bits_base_vs2_prec : _T_489;	// sequencer-master.scala:329:29
      wire [7:0] _T_554 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_522 ?
                io_op_bits_base_vs2_id : _T_490) : _T_522 ? io_op_bits_base_vs2_id : _T_490;	// sequencer-master.scala:329:29
      wire _T_555 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_523 ?
                io_op_bits_base_vs2_scalar : _T_491) : _T_523 ? io_op_bits_base_vs2_scalar : _T_491;	// sequencer-master.scala:329:29
      wire _T_556 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_524 ?
                io_op_bits_base_vs2_pred : _T_492) : _T_524 ? io_op_bits_base_vs2_pred : _T_492;	// sequencer-master.scala:329:29
      wire [1:0] _T_557 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_525 ?
                io_op_bits_base_vs2_prec : _T_493) : _T_525 ? io_op_bits_base_vs2_prec : _T_493;	// sequencer-master.scala:329:29
      wire [7:0] _T_558 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (&tail | _T_526 ?
                io_op_bits_base_vs2_id : _T_494) : _T_526 ? io_op_bits_base_vs2_id : _T_494;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_559 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (&tail | _T_527 ?
                io_op_bits_base_vs2_scalar : _T_495) : _T_527 ? io_op_bits_base_vs2_scalar : _T_495;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_560 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (&tail | _T_528 ?
                io_op_bits_base_vs2_pred : _T_496) : _T_528 ? io_op_bits_base_vs2_pred : _T_496;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_561 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid ? (&tail | _T_529 ?
                io_op_bits_base_vs2_prec : _T_497) : _T_529 ? io_op_bits_base_vs2_prec : _T_497;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_562 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_563 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_564 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_565 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_566 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_567 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_568 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_569 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_570 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_571 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_572 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_573 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_574 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_575 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_576 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_577 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_578 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_579 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_580 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_581 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_582 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_583 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_584 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_585 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_586 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_587 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_588 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_589 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_590 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_591 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_592 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_593 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_594 = (~io_op_bits_active_vint | ~_T_4) & e_0_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_595 = (~io_op_bits_active_vint | ~_T_5) & e_1_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_596 = (~io_op_bits_active_vint | ~_T_6) & e_2_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_597 = (~io_op_bits_active_vint | ~_T_7) & e_3_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_598 = (~io_op_bits_active_vint | ~_T_8) & e_4_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_599 = (~io_op_bits_active_vint | ~_T_9) & e_5_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_600 = (~io_op_bits_active_vint | ~_T_10) & e_6_base_vs3_valid;	// sequencer-master.scala:136:44, :275:29
      wire _T_601 = (~io_op_bits_active_vint | ~(&tail)) & e_7_base_vs3_valid;	// sequencer-master.scala:136:44, :267:35, :275:29, util.scala:94:11
      wire _T_602 = io_op_bits_active_vint & _T_4;	// sequencer-master.scala:289:23
      wire _T_603 = io_op_bits_active_vint & _T_5;	// sequencer-master.scala:289:23
      wire _T_604 = io_op_bits_active_vint & _T_6;	// sequencer-master.scala:289:23
      wire _T_605 = io_op_bits_active_vint & _T_7;	// sequencer-master.scala:289:23
      wire _T_606 = io_op_bits_active_vint & _T_8;	// sequencer-master.scala:289:23
      wire _T_607 = io_op_bits_active_vint & _T_9;	// sequencer-master.scala:289:23
      wire _T_608 = io_op_bits_active_vint & _T_10;	// sequencer-master.scala:289:23
      wire _T_609 = io_op_bits_active_vint & &tail;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire _T_610 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_611 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_612 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_613 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_614 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_615 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_616 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_617 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_618 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_619 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_620 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_621 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_622 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_623 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_624 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_625 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_626 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_627 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_628 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_629 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_630 = io_op_bits_active_vint & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_631 = io_op_bits_active_vint & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_632 = io_op_bits_active_vint & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_633 = io_op_bits_active_vint & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_634 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid :
                ~_T_4 & e_0_base_vs2_valid) : e_0_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_635 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid :
                ~_T_5 & e_1_base_vs2_valid) : e_1_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_636 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid :
                ~_T_6 & e_2_base_vs2_valid) : e_2_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_637 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid :
                ~_T_7 & e_3_base_vs2_valid) : e_3_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_638 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid :
                ~_T_8 & e_4_base_vs2_valid) : e_4_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_639 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid :
                ~_T_9 & e_5_base_vs2_valid) : e_5_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_640 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid :
                ~_T_10 & e_6_base_vs2_valid) : e_6_base_vs2_valid;	// sequencer-master.scala:136:44, :274:29, :329:29
      wire _T_641 = io_op_bits_active_vint ? (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid :
                ~(&tail) & e_7_base_vs2_valid) : e_7_base_vs2_valid;	// sequencer-master.scala:136:44, :267:35, :274:29, :329:29, util.scala:94:11
      wire _T_642 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_643 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & e_0_base_vd_valid) : e_0_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_644 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_645 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_646 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_647 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_648 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & e_1_base_vd_valid) : e_1_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_649 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_650 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_651 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_652 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_653 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & e_2_base_vd_valid) : e_2_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_654 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_655 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_656 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_657 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_658 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & e_3_base_vd_valid) : e_3_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_659 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_660 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_661 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_662 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_663 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & e_4_base_vd_valid) : e_4_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_664 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_665 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_666 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_667 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_668 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & e_5_base_vd_valid) : e_5_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_669 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_670 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_671 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_672 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_673 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & e_6_base_vd_valid) : e_6_base_vd_valid;	// sequencer-master.scala:136:44, :276:28, :363:24
      wire _T_674 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_675 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_676 = io_op_bits_active_vint & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_677 = io_op_bits_active_vint & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_678 = io_op_bits_active_vint ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & e_7_base_vd_valid) : e_7_base_vd_valid;	// sequencer-master.scala:136:44, :267:35, :276:28, :363:24, util.scala:94:11
      wire _T_679 = io_op_bits_active_vint & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_680 = io_op_bits_active_vint & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_681 = io_op_bits_active_vint & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_682 = (~io_op_bits_active_vipred | ~_T_4) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_4 ? io_op_bits_base_vp_valid : ~_T_4 & e_0_base_vp_valid) : e_0_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_683 = (~io_op_bits_active_vipred | ~_T_5) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_5 ? io_op_bits_base_vp_valid : ~_T_5 & e_1_base_vp_valid) : e_1_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_684 = (~io_op_bits_active_vipred | ~_T_6) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_6 ? io_op_bits_base_vp_valid : ~_T_6 & e_2_base_vp_valid) : e_2_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_685 = (~io_op_bits_active_vipred | ~_T_7) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_7 ? io_op_bits_base_vp_valid : ~_T_7 & e_3_base_vp_valid) : e_3_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_686 = (~io_op_bits_active_vipred | ~_T_8) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_8 ? io_op_bits_base_vp_valid : ~_T_8 & e_4_base_vp_valid) : e_4_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_687 = (~io_op_bits_active_vipred | ~_T_9) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid &
                _T_9 ? io_op_bits_base_vp_valid : ~_T_9 & e_5_base_vp_valid) : e_5_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_688 = (~io_op_bits_active_vipred | ~_T_10) & (io_op_bits_active_vint ? (io_op_bits_base_vp_valid
                & _T_10 ? io_op_bits_base_vp_valid : ~_T_10 & e_6_base_vp_valid) : e_6_base_vp_valid);	// sequencer-master.scala:136:44, :272:28, :321:24
      wire _T_689 = (~io_op_bits_active_vipred | ~(&tail)) & (io_op_bits_active_vint ?
                (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid : ~(&tail) &
                e_7_base_vp_valid) : e_7_base_vp_valid);	// sequencer-master.scala:136:44, :267:35, :272:28, :321:24, util.scala:94:11
      wire _T_690 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid :
                ~_T_4 & _T_634) : _T_634;	// sequencer-master.scala:274:29, :329:29
      wire _T_691 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid :
                ~_T_5 & _T_635) : _T_635;	// sequencer-master.scala:274:29, :329:29
      wire _T_692 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid :
                ~_T_6 & _T_636) : _T_636;	// sequencer-master.scala:274:29, :329:29
      wire _T_693 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid :
                ~_T_7 & _T_637) : _T_637;	// sequencer-master.scala:274:29, :329:29
      wire _T_694 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid :
                ~_T_8 & _T_638) : _T_638;	// sequencer-master.scala:274:29, :329:29
      wire _T_695 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid :
                ~_T_9 & _T_639) : _T_639;	// sequencer-master.scala:274:29, :329:29
      wire _T_696 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid :
                ~_T_10 & _T_640) : _T_640;	// sequencer-master.scala:274:29, :329:29
      wire _T_697 = io_op_bits_active_vipred ? (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid :
                ~(&tail) & _T_641) : _T_641;	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      wire [7:0] _T_698 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_4 | _T_642 ?
                io_op_bits_base_vd_id : e_0_base_vd_id) : _T_642 ? io_op_bits_base_vd_id : e_0_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_699 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & _T_643) : _T_643;	// sequencer-master.scala:276:28, :363:24
      wire _T_700 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_4 | _T_644 ?
                io_op_bits_base_vd_scalar : e_0_base_vd_scalar) : _T_644 ? io_op_bits_base_vd_scalar :
                e_0_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_701 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_4 | _T_645 ?
                io_op_bits_base_vd_pred : e_0_base_vd_pred) : _T_645 ? io_op_bits_base_vd_pred :
                e_0_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_702 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_4 | _T_646 ?
                io_op_bits_base_vd_prec : e_0_base_vd_prec) : _T_646 ? io_op_bits_base_vd_prec :
                e_0_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_703 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_5 | _T_647 ?
                io_op_bits_base_vd_id : e_1_base_vd_id) : _T_647 ? io_op_bits_base_vd_id : e_1_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_704 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & _T_648) : _T_648;	// sequencer-master.scala:276:28, :363:24
      wire _T_705 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_5 | _T_649 ?
                io_op_bits_base_vd_scalar : e_1_base_vd_scalar) : _T_649 ? io_op_bits_base_vd_scalar :
                e_1_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_706 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_5 | _T_650 ?
                io_op_bits_base_vd_pred : e_1_base_vd_pred) : _T_650 ? io_op_bits_base_vd_pred :
                e_1_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_707 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_5 | _T_651 ?
                io_op_bits_base_vd_prec : e_1_base_vd_prec) : _T_651 ? io_op_bits_base_vd_prec :
                e_1_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_708 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_6 | _T_652 ?
                io_op_bits_base_vd_id : e_2_base_vd_id) : _T_652 ? io_op_bits_base_vd_id : e_2_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_709 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & _T_653) : _T_653;	// sequencer-master.scala:276:28, :363:24
      wire _T_710 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_6 | _T_654 ?
                io_op_bits_base_vd_scalar : e_2_base_vd_scalar) : _T_654 ? io_op_bits_base_vd_scalar :
                e_2_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_711 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_6 | _T_655 ?
                io_op_bits_base_vd_pred : e_2_base_vd_pred) : _T_655 ? io_op_bits_base_vd_pred :
                e_2_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_712 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_6 | _T_656 ?
                io_op_bits_base_vd_prec : e_2_base_vd_prec) : _T_656 ? io_op_bits_base_vd_prec :
                e_2_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_713 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_7 | _T_657 ?
                io_op_bits_base_vd_id : e_3_base_vd_id) : _T_657 ? io_op_bits_base_vd_id : e_3_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_714 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & _T_658) : _T_658;	// sequencer-master.scala:276:28, :363:24
      wire _T_715 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_7 | _T_659 ?
                io_op_bits_base_vd_scalar : e_3_base_vd_scalar) : _T_659 ? io_op_bits_base_vd_scalar :
                e_3_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_716 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_7 | _T_660 ?
                io_op_bits_base_vd_pred : e_3_base_vd_pred) : _T_660 ? io_op_bits_base_vd_pred :
                e_3_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_717 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_7 | _T_661 ?
                io_op_bits_base_vd_prec : e_3_base_vd_prec) : _T_661 ? io_op_bits_base_vd_prec :
                e_3_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_718 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_8 | _T_662 ?
                io_op_bits_base_vd_id : e_4_base_vd_id) : _T_662 ? io_op_bits_base_vd_id : e_4_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_719 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & _T_663) : _T_663;	// sequencer-master.scala:276:28, :363:24
      wire _T_720 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_8 | _T_664 ?
                io_op_bits_base_vd_scalar : e_4_base_vd_scalar) : _T_664 ? io_op_bits_base_vd_scalar :
                e_4_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_721 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_8 | _T_665 ?
                io_op_bits_base_vd_pred : e_4_base_vd_pred) : _T_665 ? io_op_bits_base_vd_pred :
                e_4_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_722 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_8 | _T_666 ?
                io_op_bits_base_vd_prec : e_4_base_vd_prec) : _T_666 ? io_op_bits_base_vd_prec :
                e_4_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_723 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_9 | _T_667 ?
                io_op_bits_base_vd_id : e_5_base_vd_id) : _T_667 ? io_op_bits_base_vd_id : e_5_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_724 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & _T_668) : _T_668;	// sequencer-master.scala:276:28, :363:24
      wire _T_725 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_9 | _T_669 ?
                io_op_bits_base_vd_scalar : e_5_base_vd_scalar) : _T_669 ? io_op_bits_base_vd_scalar :
                e_5_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_726 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_9 | _T_670 ?
                io_op_bits_base_vd_pred : e_5_base_vd_pred) : _T_670 ? io_op_bits_base_vd_pred :
                e_5_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_727 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_9 | _T_671 ?
                io_op_bits_base_vd_prec : e_5_base_vd_prec) : _T_671 ? io_op_bits_base_vd_prec :
                e_5_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_728 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_10 | _T_672 ?
                io_op_bits_base_vd_id : e_6_base_vd_id) : _T_672 ? io_op_bits_base_vd_id : e_6_base_vd_id;	// sequencer-master.scala:141:29, :363:24
      wire _T_729 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & _T_673) : _T_673;	// sequencer-master.scala:276:28, :363:24
      wire _T_730 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_10 | _T_674 ?
                io_op_bits_base_vd_scalar : e_6_base_vd_scalar) : _T_674 ? io_op_bits_base_vd_scalar :
                e_6_base_vd_scalar;	// sequencer-master.scala:363:24, types-vxu.scala:119:37
      wire _T_731 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_10 | _T_675 ?
                io_op_bits_base_vd_pred : e_6_base_vd_pred) : _T_675 ? io_op_bits_base_vd_pred :
                e_6_base_vd_pred;	// sequencer-master.scala:363:24, types-vxu.scala:119:31
      wire [1:0] _T_732 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (_T_10 | _T_676 ?
                io_op_bits_base_vd_prec : e_6_base_vd_prec) : _T_676 ? io_op_bits_base_vd_prec :
                e_6_base_vd_prec;	// sequencer-master.scala:363:24
      wire [7:0] _T_733 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (&tail | _T_677 ?
                io_op_bits_base_vd_id : e_7_base_vd_id) : _T_677 ? io_op_bits_base_vd_id : e_7_base_vd_id;	// sequencer-master.scala:141:29, :267:35, :363:24, util.scala:94:11
      wire _T_734 = io_op_bits_active_vipred ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & _T_678) : _T_678;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_735 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (&tail | _T_679 ?
                io_op_bits_base_vd_scalar : e_7_base_vd_scalar) : _T_679 ? io_op_bits_base_vd_scalar :
                e_7_base_vd_scalar;	// sequencer-master.scala:267:35, :363:24, types-vxu.scala:119:37, util.scala:94:11
      wire _T_736 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (&tail | _T_680 ?
                io_op_bits_base_vd_pred : e_7_base_vd_pred) : _T_680 ? io_op_bits_base_vd_pred :
                e_7_base_vd_pred;	// sequencer-master.scala:267:35, :363:24, types-vxu.scala:119:31, util.scala:94:11
      wire [1:0] _T_737 = io_op_bits_active_vipred & io_op_bits_base_vd_valid ? (&tail | _T_681 ?
                io_op_bits_base_vd_prec : e_7_base_vd_prec) : _T_681 ? io_op_bits_base_vd_prec :
                e_7_base_vd_prec;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire [9:0] _T_738 = io_op_bits_active_vimul & _T_4 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_4 |
                _T_602 ? io_op_bits_fn_union : e_0_fn_union) : _T_602 ? io_op_bits_fn_union : e_0_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_739 = io_op_bits_active_vimul & _T_5 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_5 |
                _T_603 ? io_op_bits_fn_union : e_1_fn_union) : _T_603 ? io_op_bits_fn_union : e_1_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_740 = io_op_bits_active_vimul & _T_6 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_6 |
                _T_604 ? io_op_bits_fn_union : e_2_fn_union) : _T_604 ? io_op_bits_fn_union : e_2_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_741 = io_op_bits_active_vimul & _T_7 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_7 |
                _T_605 ? io_op_bits_fn_union : e_3_fn_union) : _T_605 ? io_op_bits_fn_union : e_3_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_742 = io_op_bits_active_vimul & _T_8 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_8 |
                _T_606 ? io_op_bits_fn_union : e_4_fn_union) : _T_606 ? io_op_bits_fn_union : e_4_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_743 = io_op_bits_active_vimul & _T_9 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_9 |
                _T_607 ? io_op_bits_fn_union : e_5_fn_union) : _T_607 ? io_op_bits_fn_union : e_5_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_744 = io_op_bits_active_vimul & _T_10 ? io_op_bits_fn_union : io_op_bits_active_vipred ? (_T_10 |
                _T_608 ? io_op_bits_fn_union : e_6_fn_union) : _T_608 ? io_op_bits_fn_union : e_6_fn_union;	// sequencer-master.scala:289:23
      wire [9:0] _T_745 = io_op_bits_active_vimul & &tail ? io_op_bits_fn_union : io_op_bits_active_vipred ? (&tail |
                _T_609 ? io_op_bits_fn_union : e_7_fn_union) : _T_609 ? io_op_bits_fn_union : e_7_fn_union;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire [3:0] _T_746 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_4 | _T_610 ? io_op_bits_base_vp_id
                : e_0_base_vp_id) : _T_610 ? io_op_bits_base_vp_id : e_0_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_747 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_682) : _T_682;	// sequencer-master.scala:272:28, :321:24
      wire _T_748 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_4 | _T_611 ?
                io_op_bits_base_vp_scalar : e_0_base_vp_scalar) : _T_611 ? io_op_bits_base_vp_scalar :
                e_0_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_749 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_4 | _T_612 ?
                io_op_bits_base_vp_pred : e_0_base_vp_pred) : _T_612 ? io_op_bits_base_vp_pred :
                e_0_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_750 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_5 | _T_613 ? io_op_bits_base_vp_id
                : e_1_base_vp_id) : _T_613 ? io_op_bits_base_vp_id : e_1_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_751 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_683) : _T_683;	// sequencer-master.scala:272:28, :321:24
      wire _T_752 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_5 | _T_614 ?
                io_op_bits_base_vp_scalar : e_1_base_vp_scalar) : _T_614 ? io_op_bits_base_vp_scalar :
                e_1_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_753 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_5 | _T_615 ?
                io_op_bits_base_vp_pred : e_1_base_vp_pred) : _T_615 ? io_op_bits_base_vp_pred :
                e_1_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_754 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_6 | _T_616 ? io_op_bits_base_vp_id
                : e_2_base_vp_id) : _T_616 ? io_op_bits_base_vp_id : e_2_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_755 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_684) : _T_684;	// sequencer-master.scala:272:28, :321:24
      wire _T_756 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_6 | _T_617 ?
                io_op_bits_base_vp_scalar : e_2_base_vp_scalar) : _T_617 ? io_op_bits_base_vp_scalar :
                e_2_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_757 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_6 | _T_618 ?
                io_op_bits_base_vp_pred : e_2_base_vp_pred) : _T_618 ? io_op_bits_base_vp_pred :
                e_2_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_758 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_7 | _T_619 ? io_op_bits_base_vp_id
                : e_3_base_vp_id) : _T_619 ? io_op_bits_base_vp_id : e_3_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_759 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_685) : _T_685;	// sequencer-master.scala:272:28, :321:24
      wire _T_760 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_7 | _T_620 ?
                io_op_bits_base_vp_scalar : e_3_base_vp_scalar) : _T_620 ? io_op_bits_base_vp_scalar :
                e_3_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_761 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_7 | _T_621 ?
                io_op_bits_base_vp_pred : e_3_base_vp_pred) : _T_621 ? io_op_bits_base_vp_pred :
                e_3_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_762 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_8 | _T_622 ? io_op_bits_base_vp_id
                : e_4_base_vp_id) : _T_622 ? io_op_bits_base_vp_id : e_4_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_763 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_686) : _T_686;	// sequencer-master.scala:272:28, :321:24
      wire _T_764 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_8 | _T_623 ?
                io_op_bits_base_vp_scalar : e_4_base_vp_scalar) : _T_623 ? io_op_bits_base_vp_scalar :
                e_4_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_765 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_8 | _T_624 ?
                io_op_bits_base_vp_pred : e_4_base_vp_pred) : _T_624 ? io_op_bits_base_vp_pred :
                e_4_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_766 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_9 | _T_625 ? io_op_bits_base_vp_id
                : e_5_base_vp_id) : _T_625 ? io_op_bits_base_vp_id : e_5_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_767 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_687) : _T_687;	// sequencer-master.scala:272:28, :321:24
      wire _T_768 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_9 | _T_626 ?
                io_op_bits_base_vp_scalar : e_5_base_vp_scalar) : _T_626 ? io_op_bits_base_vp_scalar :
                e_5_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_769 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_9 | _T_627 ?
                io_op_bits_base_vp_pred : e_5_base_vp_pred) : _T_627 ? io_op_bits_base_vp_pred :
                e_5_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_770 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_10 | _T_628 ?
                io_op_bits_base_vp_id : e_6_base_vp_id) : _T_628 ? io_op_bits_base_vp_id : e_6_base_vp_id;	// sequencer-master.scala:141:29, :321:24
      wire _T_771 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_688) : _T_688;	// sequencer-master.scala:272:28, :321:24
      wire _T_772 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_10 | _T_629 ?
                io_op_bits_base_vp_scalar : e_6_base_vp_scalar) : _T_629 ? io_op_bits_base_vp_scalar :
                e_6_base_vp_scalar;	// sequencer-master.scala:321:24, types-vxu.scala:119:37
      wire _T_773 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (_T_10 | _T_630 ?
                io_op_bits_base_vp_pred : e_6_base_vp_pred) : _T_630 ? io_op_bits_base_vp_pred :
                e_6_base_vp_pred;	// sequencer-master.scala:321:24, types-vxu.scala:119:31
      wire [3:0] _T_774 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (&tail | _T_631 ?
                io_op_bits_base_vp_id : e_7_base_vp_id) : _T_631 ? io_op_bits_base_vp_id : e_7_base_vp_id;	// sequencer-master.scala:141:29, :267:35, :321:24, util.scala:94:11
      wire _T_775 = io_op_bits_active_vimul ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_689) : _T_689;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_776 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (&tail | _T_632 ?
                io_op_bits_base_vp_scalar : e_7_base_vp_scalar) : _T_632 ? io_op_bits_base_vp_scalar :
                e_7_base_vp_scalar;	// sequencer-master.scala:267:35, :321:24, types-vxu.scala:119:37, util.scala:94:11
      wire _T_777 = io_op_bits_active_vimul & io_op_bits_base_vp_valid ? (&tail | _T_633 ?
                io_op_bits_base_vp_pred : e_7_base_vp_pred) : _T_633 ? io_op_bits_base_vp_pred :
                e_7_base_vp_pred;	// sequencer-master.scala:267:35, :321:24, types-vxu.scala:119:31, util.scala:94:11
      wire _T_778 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid :
                ~_T_4 & _T_690) : _T_690;	// sequencer-master.scala:274:29, :329:29
      wire _T_779 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid :
                ~_T_5 & _T_691) : _T_691;	// sequencer-master.scala:274:29, :329:29
      wire _T_780 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid :
                ~_T_6 & _T_692) : _T_692;	// sequencer-master.scala:274:29, :329:29
      wire _T_781 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid :
                ~_T_7 & _T_693) : _T_693;	// sequencer-master.scala:274:29, :329:29
      wire _T_782 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid :
                ~_T_8 & _T_694) : _T_694;	// sequencer-master.scala:274:29, :329:29
      wire _T_783 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid :
                ~_T_9 & _T_695) : _T_695;	// sequencer-master.scala:274:29, :329:29
      wire _T_784 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid :
                ~_T_10 & _T_696) : _T_696;	// sequencer-master.scala:274:29, :329:29
      wire _T_785 = io_op_bits_active_vimul ? (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid :
                ~(&tail) & _T_697) : _T_697;	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      wire _T_786 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_787 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & _T_699) : _T_699;	// sequencer-master.scala:276:28, :363:24
      wire _T_788 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_789 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_790 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_791 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_792 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & _T_704) : _T_704;	// sequencer-master.scala:276:28, :363:24
      wire _T_793 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_794 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_795 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_796 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_797 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & _T_709) : _T_709;	// sequencer-master.scala:276:28, :363:24
      wire _T_798 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_799 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_800 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_801 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_802 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & _T_714) : _T_714;	// sequencer-master.scala:276:28, :363:24
      wire _T_803 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_804 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_805 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_806 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_807 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & _T_719) : _T_719;	// sequencer-master.scala:276:28, :363:24
      wire _T_808 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_809 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_810 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_811 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_812 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & _T_724) : _T_724;	// sequencer-master.scala:276:28, :363:24
      wire _T_813 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_814 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_815 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_816 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_817 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & _T_729) : _T_729;	// sequencer-master.scala:276:28, :363:24
      wire _T_818 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_819 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_820 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_821 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_822 = io_op_bits_active_vimul ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & _T_734) : _T_734;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_823 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_824 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_825 = io_op_bits_active_vimul & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_826 = _T_107 | io_op_bits_active_vrfirst;	// sequencer-master.scala:301:46
      wire [9:0] _T_827 = {8'h0, io_op_bits_active_vidiv | io_op_bits_active_vfdiv & ~(io_op_bits_fn_union[0]),
                _T_826};	// sequencer-master.scala:289:23, :300:{28,46}, :411:70, types-vxu.scala:54:51, :96:47
      wire _T_828 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_829 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_830 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_831 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_832 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_833 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_834 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_835 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_836 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_837 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_838 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_839 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_840 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_841 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_842 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_843 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_844 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_845 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_846 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_847 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_848 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_849 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_850 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_851 = io_op_bits_active_vidiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_852 = io_op_bits_active_vidiv ? ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ?
                io_op_bits_base_vp_valid : ~_T_4 & _T_747) : _T_747;	// sequencer-master.scala:272:28, :321:24
      wire _T_853 = io_op_bits_active_vidiv ? ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ?
                io_op_bits_base_vp_valid : ~_T_5 & _T_751) : _T_751;	// sequencer-master.scala:272:28, :321:24
      wire _T_854 = io_op_bits_active_vidiv ? ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ?
                io_op_bits_base_vp_valid : ~_T_6 & _T_755) : _T_755;	// sequencer-master.scala:272:28, :321:24
      wire _T_855 = io_op_bits_active_vidiv ? ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ?
                io_op_bits_base_vp_valid : ~_T_7 & _T_759) : _T_759;	// sequencer-master.scala:272:28, :321:24
      wire _T_856 = io_op_bits_active_vidiv ? ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ?
                io_op_bits_base_vp_valid : ~_T_8 & _T_763) : _T_763;	// sequencer-master.scala:272:28, :321:24
      wire _T_857 = io_op_bits_active_vidiv ? ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ?
                io_op_bits_base_vp_valid : ~_T_9 & _T_767) : _T_767;	// sequencer-master.scala:272:28, :321:24
      wire _T_858 = io_op_bits_active_vidiv ? ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ?
                io_op_bits_base_vp_valid : ~_T_10 & _T_771) : _T_771;	// sequencer-master.scala:272:28, :321:24
      wire _T_859 = io_op_bits_active_vidiv ? ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ?
                io_op_bits_base_vp_valid : ~(&tail) & _T_775) : _T_775;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_860 = io_op_bits_active_vidiv ? ~_T_132 & (io_op_bits_base_vs2_valid & _T_4 ?
                io_op_bits_base_vs2_valid : ~_T_4 & _T_778) : _T_778;	// sequencer-master.scala:274:29, :329:29
      wire _T_861 = io_op_bits_active_vidiv ? ~_T_133 & (io_op_bits_base_vs2_valid & _T_5 ?
                io_op_bits_base_vs2_valid : ~_T_5 & _T_779) : _T_779;	// sequencer-master.scala:274:29, :329:29
      wire _T_862 = io_op_bits_active_vidiv ? ~_T_134 & (io_op_bits_base_vs2_valid & _T_6 ?
                io_op_bits_base_vs2_valid : ~_T_6 & _T_780) : _T_780;	// sequencer-master.scala:274:29, :329:29
      wire _T_863 = io_op_bits_active_vidiv ? ~_T_135 & (io_op_bits_base_vs2_valid & _T_7 ?
                io_op_bits_base_vs2_valid : ~_T_7 & _T_781) : _T_781;	// sequencer-master.scala:274:29, :329:29
      wire _T_864 = io_op_bits_active_vidiv ? ~_T_136 & (io_op_bits_base_vs2_valid & _T_8 ?
                io_op_bits_base_vs2_valid : ~_T_8 & _T_782) : _T_782;	// sequencer-master.scala:274:29, :329:29
      wire _T_865 = io_op_bits_active_vidiv ? ~_T_137 & (io_op_bits_base_vs2_valid & _T_9 ?
                io_op_bits_base_vs2_valid : ~_T_9 & _T_783) : _T_783;	// sequencer-master.scala:274:29, :329:29
      wire _T_866 = io_op_bits_active_vidiv ? ~_T_138 & (io_op_bits_base_vs2_valid & _T_10 ?
                io_op_bits_base_vs2_valid : ~_T_10 & _T_784) : _T_784;	// sequencer-master.scala:274:29, :329:29
      wire _T_867 = io_op_bits_active_vidiv ? ~(&_T_0) & (io_op_bits_base_vs2_valid & &tail ?
                io_op_bits_base_vs2_valid : ~(&tail) & _T_785) : _T_785;	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      wire _T_868 = (~io_op_bits_active_vidiv | ~_T_132 & ~_T_4) & (~io_op_bits_active_vimul | ~_T_4) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_4 ? io_op_bits_base_vs3_valid :
                ~_T_4 & _T_594) : _T_594);	// sequencer-master.scala:275:29, :329:29
      wire _T_869 = (~io_op_bits_active_vidiv | ~_T_133 & ~_T_5) & (~io_op_bits_active_vimul | ~_T_5) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_5 ? io_op_bits_base_vs3_valid :
                ~_T_5 & _T_595) : _T_595);	// sequencer-master.scala:275:29, :329:29
      wire _T_870 = (~io_op_bits_active_vidiv | ~_T_134 & ~_T_6) & (~io_op_bits_active_vimul | ~_T_6) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_6 ? io_op_bits_base_vs3_valid :
                ~_T_6 & _T_596) : _T_596);	// sequencer-master.scala:275:29, :329:29
      wire _T_871 = (~io_op_bits_active_vidiv | ~_T_135 & ~_T_7) & (~io_op_bits_active_vimul | ~_T_7) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_7 ? io_op_bits_base_vs3_valid :
                ~_T_7 & _T_597) : _T_597);	// sequencer-master.scala:275:29, :329:29
      wire _T_872 = (~io_op_bits_active_vidiv | ~_T_136 & ~_T_8) & (~io_op_bits_active_vimul | ~_T_8) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_8 ? io_op_bits_base_vs3_valid :
                ~_T_8 & _T_598) : _T_598);	// sequencer-master.scala:275:29, :329:29
      wire _T_873 = (~io_op_bits_active_vidiv | ~_T_137 & ~_T_9) & (~io_op_bits_active_vimul | ~_T_9) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_9 ? io_op_bits_base_vs3_valid :
                ~_T_9 & _T_599) : _T_599);	// sequencer-master.scala:275:29, :329:29
      wire _T_874 = (~io_op_bits_active_vidiv | ~_T_138 & ~_T_10) & (~io_op_bits_active_vimul | ~_T_10) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & _T_10 ? io_op_bits_base_vs3_valid
                : ~_T_10 & _T_600) : _T_600);	// sequencer-master.scala:275:29, :329:29
      wire _T_875 = (~io_op_bits_active_vidiv | ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vimul | ~(&tail)) &
                (io_op_bits_active_vipred ? (io_op_bits_base_vs3_valid & &tail ? io_op_bits_base_vs3_valid
                : ~(&tail) & _T_601) : _T_601);	// sequencer-master.scala:267:35, :275:29, :329:29, util.scala:94:11
      wire [7:0] _T_876 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_132 | _T_786 ?
                io_op_bits_base_vd_id : _T_698) : _T_786 ? io_op_bits_base_vd_id : _T_698;	// sequencer-master.scala:363:24
      wire _T_877 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_132 ? io_op_bits_base_vd_valid :
                ~_T_132 & ~_T_4 & _T_787) : _T_787;	// sequencer-master.scala:276:28, :363:24
      wire _T_878 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_132 | _T_788 ?
                io_op_bits_base_vd_scalar : _T_700) : _T_788 ? io_op_bits_base_vd_scalar : _T_700;	// sequencer-master.scala:363:24
      wire _T_879 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_132 | _T_789 ?
                io_op_bits_base_vd_pred : _T_701) : _T_789 ? io_op_bits_base_vd_pred : _T_701;	// sequencer-master.scala:363:24
      wire [1:0] _T_880 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_132 | _T_790 ?
                io_op_bits_base_vd_prec : _T_702) : _T_790 ? io_op_bits_base_vd_prec : _T_702;	// sequencer-master.scala:363:24
      wire [7:0] _T_881 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_133 | _T_791 ?
                io_op_bits_base_vd_id : _T_703) : _T_791 ? io_op_bits_base_vd_id : _T_703;	// sequencer-master.scala:363:24
      wire _T_882 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_133 ? io_op_bits_base_vd_valid :
                ~_T_133 & ~_T_5 & _T_792) : _T_792;	// sequencer-master.scala:276:28, :363:24
      wire _T_883 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_133 | _T_793 ?
                io_op_bits_base_vd_scalar : _T_705) : _T_793 ? io_op_bits_base_vd_scalar : _T_705;	// sequencer-master.scala:363:24
      wire _T_884 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_133 | _T_794 ?
                io_op_bits_base_vd_pred : _T_706) : _T_794 ? io_op_bits_base_vd_pred : _T_706;	// sequencer-master.scala:363:24
      wire [1:0] _T_885 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_133 | _T_795 ?
                io_op_bits_base_vd_prec : _T_707) : _T_795 ? io_op_bits_base_vd_prec : _T_707;	// sequencer-master.scala:363:24
      wire [7:0] _T_886 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_134 | _T_796 ?
                io_op_bits_base_vd_id : _T_708) : _T_796 ? io_op_bits_base_vd_id : _T_708;	// sequencer-master.scala:363:24
      wire _T_887 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_134 ? io_op_bits_base_vd_valid :
                ~_T_134 & ~_T_6 & _T_797) : _T_797;	// sequencer-master.scala:276:28, :363:24
      wire _T_888 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_134 | _T_798 ?
                io_op_bits_base_vd_scalar : _T_710) : _T_798 ? io_op_bits_base_vd_scalar : _T_710;	// sequencer-master.scala:363:24
      wire _T_889 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_134 | _T_799 ?
                io_op_bits_base_vd_pred : _T_711) : _T_799 ? io_op_bits_base_vd_pred : _T_711;	// sequencer-master.scala:363:24
      wire [1:0] _T_890 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_134 | _T_800 ?
                io_op_bits_base_vd_prec : _T_712) : _T_800 ? io_op_bits_base_vd_prec : _T_712;	// sequencer-master.scala:363:24
      wire [7:0] _T_891 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_135 | _T_801 ?
                io_op_bits_base_vd_id : _T_713) : _T_801 ? io_op_bits_base_vd_id : _T_713;	// sequencer-master.scala:363:24
      wire _T_892 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_135 ? io_op_bits_base_vd_valid :
                ~_T_135 & ~_T_7 & _T_802) : _T_802;	// sequencer-master.scala:276:28, :363:24
      wire _T_893 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_135 | _T_803 ?
                io_op_bits_base_vd_scalar : _T_715) : _T_803 ? io_op_bits_base_vd_scalar : _T_715;	// sequencer-master.scala:363:24
      wire _T_894 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_135 | _T_804 ?
                io_op_bits_base_vd_pred : _T_716) : _T_804 ? io_op_bits_base_vd_pred : _T_716;	// sequencer-master.scala:363:24
      wire [1:0] _T_895 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_135 | _T_805 ?
                io_op_bits_base_vd_prec : _T_717) : _T_805 ? io_op_bits_base_vd_prec : _T_717;	// sequencer-master.scala:363:24
      wire [7:0] _T_896 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_136 | _T_806 ?
                io_op_bits_base_vd_id : _T_718) : _T_806 ? io_op_bits_base_vd_id : _T_718;	// sequencer-master.scala:363:24
      wire _T_897 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_136 ? io_op_bits_base_vd_valid :
                ~_T_136 & ~_T_8 & _T_807) : _T_807;	// sequencer-master.scala:276:28, :363:24
      wire _T_898 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_136 | _T_808 ?
                io_op_bits_base_vd_scalar : _T_720) : _T_808 ? io_op_bits_base_vd_scalar : _T_720;	// sequencer-master.scala:363:24
      wire _T_899 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_136 | _T_809 ?
                io_op_bits_base_vd_pred : _T_721) : _T_809 ? io_op_bits_base_vd_pred : _T_721;	// sequencer-master.scala:363:24
      wire [1:0] _T_900 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_136 | _T_810 ?
                io_op_bits_base_vd_prec : _T_722) : _T_810 ? io_op_bits_base_vd_prec : _T_722;	// sequencer-master.scala:363:24
      wire [7:0] _T_901 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_137 | _T_811 ?
                io_op_bits_base_vd_id : _T_723) : _T_811 ? io_op_bits_base_vd_id : _T_723;	// sequencer-master.scala:363:24
      wire _T_902 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_137 ? io_op_bits_base_vd_valid :
                ~_T_137 & ~_T_9 & _T_812) : _T_812;	// sequencer-master.scala:276:28, :363:24
      wire _T_903 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_137 | _T_813 ?
                io_op_bits_base_vd_scalar : _T_725) : _T_813 ? io_op_bits_base_vd_scalar : _T_725;	// sequencer-master.scala:363:24
      wire _T_904 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_137 | _T_814 ?
                io_op_bits_base_vd_pred : _T_726) : _T_814 ? io_op_bits_base_vd_pred : _T_726;	// sequencer-master.scala:363:24
      wire [1:0] _T_905 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_137 | _T_815 ?
                io_op_bits_base_vd_prec : _T_727) : _T_815 ? io_op_bits_base_vd_prec : _T_727;	// sequencer-master.scala:363:24
      wire [7:0] _T_906 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_138 | _T_816 ?
                io_op_bits_base_vd_id : _T_728) : _T_816 ? io_op_bits_base_vd_id : _T_728;	// sequencer-master.scala:363:24
      wire _T_907 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & _T_138 ? io_op_bits_base_vd_valid :
                ~_T_138 & ~_T_10 & _T_817) : _T_817;	// sequencer-master.scala:276:28, :363:24
      wire _T_908 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_138 | _T_818 ?
                io_op_bits_base_vd_scalar : _T_730) : _T_818 ? io_op_bits_base_vd_scalar : _T_730;	// sequencer-master.scala:363:24
      wire _T_909 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_138 | _T_819 ?
                io_op_bits_base_vd_pred : _T_731) : _T_819 ? io_op_bits_base_vd_pred : _T_731;	// sequencer-master.scala:363:24
      wire [1:0] _T_910 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (_T_138 | _T_820 ?
                io_op_bits_base_vd_prec : _T_732) : _T_820 ? io_op_bits_base_vd_prec : _T_732;	// sequencer-master.scala:363:24
      wire [7:0] _T_911 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_821 ?
                io_op_bits_base_vd_id : _T_733) : _T_821 ? io_op_bits_base_vd_id : _T_733;	// sequencer-master.scala:267:35, :363:24
      wire _T_912 = io_op_bits_active_vidiv ? (io_op_bits_base_vd_valid & &_T_0 ? io_op_bits_base_vd_valid :
                ~(&_T_0) & ~(&tail) & _T_822) : _T_822;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_913 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_823 ?
                io_op_bits_base_vd_scalar : _T_735) : _T_823 ? io_op_bits_base_vd_scalar : _T_735;	// sequencer-master.scala:267:35, :363:24
      wire _T_914 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_824 ?
                io_op_bits_base_vd_pred : _T_736) : _T_824 ? io_op_bits_base_vd_pred : _T_736;	// sequencer-master.scala:267:35, :363:24
      wire [1:0] _T_915 = io_op_bits_active_vidiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_825 ?
                io_op_bits_base_vd_prec : _T_737) : _T_825 ? io_op_bits_base_vd_prec : _T_737;	// sequencer-master.scala:267:35, :363:24
      wire [9:0] _T_916 = io_op_bits_active_vfma & _T_4 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_132 ?
                io_op_bits_fn_union : _T_4 ? _T_827 : _T_738) : _T_738;	// sequencer-master.scala:289:23
      wire [9:0] _T_917 = io_op_bits_active_vfma & _T_5 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_133 ?
                io_op_bits_fn_union : _T_5 ? _T_827 : _T_739) : _T_739;	// sequencer-master.scala:289:23
      wire [9:0] _T_918 = io_op_bits_active_vfma & _T_6 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_134 ?
                io_op_bits_fn_union : _T_6 ? _T_827 : _T_740) : _T_740;	// sequencer-master.scala:289:23
      wire [9:0] _T_919 = io_op_bits_active_vfma & _T_7 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_135 ?
                io_op_bits_fn_union : _T_7 ? _T_827 : _T_741) : _T_741;	// sequencer-master.scala:289:23
      wire [9:0] _T_920 = io_op_bits_active_vfma & _T_8 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_136 ?
                io_op_bits_fn_union : _T_8 ? _T_827 : _T_742) : _T_742;	// sequencer-master.scala:289:23
      wire [9:0] _T_921 = io_op_bits_active_vfma & _T_9 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_137 ?
                io_op_bits_fn_union : _T_9 ? _T_827 : _T_743) : _T_743;	// sequencer-master.scala:289:23
      wire [9:0] _T_922 = io_op_bits_active_vfma & _T_10 ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (_T_138 ?
                io_op_bits_fn_union : _T_10 ? _T_827 : _T_744) : _T_744;	// sequencer-master.scala:289:23
      wire [9:0] _T_923 = io_op_bits_active_vfma & &tail ? io_op_bits_fn_union : io_op_bits_active_vidiv ? (&_T_0 ?
                io_op_bits_fn_union : &tail ? _T_827 : _T_745) : _T_745;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire [3:0] _T_924 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_4 | _T_828 ? io_op_bits_base_vp_id
                : _T_746) : _T_828 ? io_op_bits_base_vp_id : _T_746;	// sequencer-master.scala:321:24
      wire _T_925 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_852) : _T_852;	// sequencer-master.scala:272:28, :321:24
      wire _T_926 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_4 | _T_829 ?
                io_op_bits_base_vp_scalar : _T_748) : _T_829 ? io_op_bits_base_vp_scalar : _T_748;	// sequencer-master.scala:321:24
      wire _T_927 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_4 | _T_830 ?
                io_op_bits_base_vp_pred : _T_749) : _T_830 ? io_op_bits_base_vp_pred : _T_749;	// sequencer-master.scala:321:24
      wire [3:0] _T_928 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_5 | _T_831 ? io_op_bits_base_vp_id
                : _T_750) : _T_831 ? io_op_bits_base_vp_id : _T_750;	// sequencer-master.scala:321:24
      wire _T_929 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_853) : _T_853;	// sequencer-master.scala:272:28, :321:24
      wire _T_930 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_5 | _T_832 ?
                io_op_bits_base_vp_scalar : _T_752) : _T_832 ? io_op_bits_base_vp_scalar : _T_752;	// sequencer-master.scala:321:24
      wire _T_931 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_5 | _T_833 ?
                io_op_bits_base_vp_pred : _T_753) : _T_833 ? io_op_bits_base_vp_pred : _T_753;	// sequencer-master.scala:321:24
      wire [3:0] _T_932 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_6 | _T_834 ? io_op_bits_base_vp_id
                : _T_754) : _T_834 ? io_op_bits_base_vp_id : _T_754;	// sequencer-master.scala:321:24
      wire _T_933 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_854) : _T_854;	// sequencer-master.scala:272:28, :321:24
      wire _T_934 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_6 | _T_835 ?
                io_op_bits_base_vp_scalar : _T_756) : _T_835 ? io_op_bits_base_vp_scalar : _T_756;	// sequencer-master.scala:321:24
      wire _T_935 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_6 | _T_836 ?
                io_op_bits_base_vp_pred : _T_757) : _T_836 ? io_op_bits_base_vp_pred : _T_757;	// sequencer-master.scala:321:24
      wire [3:0] _T_936 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_7 | _T_837 ? io_op_bits_base_vp_id
                : _T_758) : _T_837 ? io_op_bits_base_vp_id : _T_758;	// sequencer-master.scala:321:24
      wire _T_937 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_855) : _T_855;	// sequencer-master.scala:272:28, :321:24
      wire _T_938 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_7 | _T_838 ?
                io_op_bits_base_vp_scalar : _T_760) : _T_838 ? io_op_bits_base_vp_scalar : _T_760;	// sequencer-master.scala:321:24
      wire _T_939 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_7 | _T_839 ?
                io_op_bits_base_vp_pred : _T_761) : _T_839 ? io_op_bits_base_vp_pred : _T_761;	// sequencer-master.scala:321:24
      wire [3:0] _T_940 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_8 | _T_840 ? io_op_bits_base_vp_id
                : _T_762) : _T_840 ? io_op_bits_base_vp_id : _T_762;	// sequencer-master.scala:321:24
      wire _T_941 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_856) : _T_856;	// sequencer-master.scala:272:28, :321:24
      wire _T_942 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_8 | _T_841 ?
                io_op_bits_base_vp_scalar : _T_764) : _T_841 ? io_op_bits_base_vp_scalar : _T_764;	// sequencer-master.scala:321:24
      wire _T_943 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_8 | _T_842 ?
                io_op_bits_base_vp_pred : _T_765) : _T_842 ? io_op_bits_base_vp_pred : _T_765;	// sequencer-master.scala:321:24
      wire [3:0] _T_944 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_9 | _T_843 ? io_op_bits_base_vp_id
                : _T_766) : _T_843 ? io_op_bits_base_vp_id : _T_766;	// sequencer-master.scala:321:24
      wire _T_945 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_857) : _T_857;	// sequencer-master.scala:272:28, :321:24
      wire _T_946 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_9 | _T_844 ?
                io_op_bits_base_vp_scalar : _T_768) : _T_844 ? io_op_bits_base_vp_scalar : _T_768;	// sequencer-master.scala:321:24
      wire _T_947 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_9 | _T_845 ?
                io_op_bits_base_vp_pred : _T_769) : _T_845 ? io_op_bits_base_vp_pred : _T_769;	// sequencer-master.scala:321:24
      wire [3:0] _T_948 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_10 | _T_846 ? io_op_bits_base_vp_id
                : _T_770) : _T_846 ? io_op_bits_base_vp_id : _T_770;	// sequencer-master.scala:321:24
      wire _T_949 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_858) : _T_858;	// sequencer-master.scala:272:28, :321:24
      wire _T_950 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_10 | _T_847 ?
                io_op_bits_base_vp_scalar : _T_772) : _T_847 ? io_op_bits_base_vp_scalar : _T_772;	// sequencer-master.scala:321:24
      wire _T_951 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (_T_10 | _T_848 ?
                io_op_bits_base_vp_pred : _T_773) : _T_848 ? io_op_bits_base_vp_pred : _T_773;	// sequencer-master.scala:321:24
      wire [3:0] _T_952 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (&tail | _T_849 ? io_op_bits_base_vp_id
                : _T_774) : _T_849 ? io_op_bits_base_vp_id : _T_774;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_953 = io_op_bits_active_vfma ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_859) : _T_859;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_954 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (&tail | _T_850 ?
                io_op_bits_base_vp_scalar : _T_776) : _T_850 ? io_op_bits_base_vp_scalar : _T_776;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_955 = io_op_bits_active_vfma & io_op_bits_base_vp_valid ? (&tail | _T_851 ?
                io_op_bits_base_vp_pred : _T_777) : _T_851 ? io_op_bits_base_vp_pred : _T_777;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_956 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid :
                ~_T_4 & _T_860) : _T_860;	// sequencer-master.scala:274:29, :329:29
      wire _T_957 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid :
                ~_T_5 & _T_861) : _T_861;	// sequencer-master.scala:274:29, :329:29
      wire _T_958 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid :
                ~_T_6 & _T_862) : _T_862;	// sequencer-master.scala:274:29, :329:29
      wire _T_959 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid :
                ~_T_7 & _T_863) : _T_863;	// sequencer-master.scala:274:29, :329:29
      wire _T_960 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid :
                ~_T_8 & _T_864) : _T_864;	// sequencer-master.scala:274:29, :329:29
      wire _T_961 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid :
                ~_T_9 & _T_865) : _T_865;	// sequencer-master.scala:274:29, :329:29
      wire _T_962 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid :
                ~_T_10 & _T_866) : _T_866;	// sequencer-master.scala:274:29, :329:29
      wire _T_963 = io_op_bits_active_vfma ? (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid :
                ~(&tail) & _T_867) : _T_867;	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      wire _T_964 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_965 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & _T_877) : _T_877;	// sequencer-master.scala:276:28, :363:24
      wire _T_966 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_967 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_968 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_969 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_970 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & _T_882) : _T_882;	// sequencer-master.scala:276:28, :363:24
      wire _T_971 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_972 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_973 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_974 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_975 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & _T_887) : _T_887;	// sequencer-master.scala:276:28, :363:24
      wire _T_976 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_977 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_978 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_979 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_980 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & _T_892) : _T_892;	// sequencer-master.scala:276:28, :363:24
      wire _T_981 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_982 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_983 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_984 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_985 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & _T_897) : _T_897;	// sequencer-master.scala:276:28, :363:24
      wire _T_986 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_987 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_988 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_989 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_990 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & _T_902) : _T_902;	// sequencer-master.scala:276:28, :363:24
      wire _T_991 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_992 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_993 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_994 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_995 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & _T_907) : _T_907;	// sequencer-master.scala:276:28, :363:24
      wire _T_996 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_997 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_998 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_999 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1000 = io_op_bits_active_vfma ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & _T_912) : _T_912;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_1001 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1002 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1003 = io_op_bits_active_vfma & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire [9:0] _T_1004 = {8'h0, io_op_bits_active_vidiv | io_op_bits_active_vfdiv & ~(io_op_bits_fn_union[0]),
                _T_826};	// sequencer-master.scala:289:23, :300:{28,46}, :411:70, types-vxu.scala:54:51, :96:47
      wire _T_1005 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1006 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1007 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1008 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1009 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1010 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1011 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1012 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1013 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1014 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1015 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1016 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1017 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1018 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1019 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1020 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1021 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1022 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1023 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1024 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1025 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1026 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1027 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1028 = io_op_bits_active_vfdiv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1029 = io_op_bits_active_vfdiv ? ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ?
                io_op_bits_base_vp_valid : ~_T_4 & _T_925) : _T_925;	// sequencer-master.scala:272:28, :321:24
      wire _T_1030 = io_op_bits_active_vfdiv ? ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ?
                io_op_bits_base_vp_valid : ~_T_5 & _T_929) : _T_929;	// sequencer-master.scala:272:28, :321:24
      wire _T_1031 = io_op_bits_active_vfdiv ? ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ?
                io_op_bits_base_vp_valid : ~_T_6 & _T_933) : _T_933;	// sequencer-master.scala:272:28, :321:24
      wire _T_1032 = io_op_bits_active_vfdiv ? ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ?
                io_op_bits_base_vp_valid : ~_T_7 & _T_937) : _T_937;	// sequencer-master.scala:272:28, :321:24
      wire _T_1033 = io_op_bits_active_vfdiv ? ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ?
                io_op_bits_base_vp_valid : ~_T_8 & _T_941) : _T_941;	// sequencer-master.scala:272:28, :321:24
      wire _T_1034 = io_op_bits_active_vfdiv ? ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ?
                io_op_bits_base_vp_valid : ~_T_9 & _T_945) : _T_945;	// sequencer-master.scala:272:28, :321:24
      wire _T_1035 = io_op_bits_active_vfdiv ? ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ?
                io_op_bits_base_vp_valid : ~_T_10 & _T_949) : _T_949;	// sequencer-master.scala:272:28, :321:24
      wire _T_1036 = io_op_bits_active_vfdiv ? ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ?
                io_op_bits_base_vp_valid : ~(&tail) & _T_953) : _T_953;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1037 = io_op_bits_active_vfdiv ? ~_T_132 & (io_op_bits_base_vs2_valid & _T_4 ?
                io_op_bits_base_vs2_valid : ~_T_4 & _T_956) : _T_956;	// sequencer-master.scala:274:29, :329:29
      wire _T_1038 = io_op_bits_active_vfdiv ? ~_T_133 & (io_op_bits_base_vs2_valid & _T_5 ?
                io_op_bits_base_vs2_valid : ~_T_5 & _T_957) : _T_957;	// sequencer-master.scala:274:29, :329:29
      wire _T_1039 = io_op_bits_active_vfdiv ? ~_T_134 & (io_op_bits_base_vs2_valid & _T_6 ?
                io_op_bits_base_vs2_valid : ~_T_6 & _T_958) : _T_958;	// sequencer-master.scala:274:29, :329:29
      wire _T_1040 = io_op_bits_active_vfdiv ? ~_T_135 & (io_op_bits_base_vs2_valid & _T_7 ?
                io_op_bits_base_vs2_valid : ~_T_7 & _T_959) : _T_959;	// sequencer-master.scala:274:29, :329:29
      wire _T_1041 = io_op_bits_active_vfdiv ? ~_T_136 & (io_op_bits_base_vs2_valid & _T_8 ?
                io_op_bits_base_vs2_valid : ~_T_8 & _T_960) : _T_960;	// sequencer-master.scala:274:29, :329:29
      wire _T_1042 = io_op_bits_active_vfdiv ? ~_T_137 & (io_op_bits_base_vs2_valid & _T_9 ?
                io_op_bits_base_vs2_valid : ~_T_9 & _T_961) : _T_961;	// sequencer-master.scala:274:29, :329:29
      wire _T_1043 = io_op_bits_active_vfdiv ? ~_T_138 & (io_op_bits_base_vs2_valid & _T_10 ?
                io_op_bits_base_vs2_valid : ~_T_10 & _T_962) : _T_962;	// sequencer-master.scala:274:29, :329:29
      wire _T_1044 = io_op_bits_active_vfdiv ? ~(&_T_0) & (io_op_bits_base_vs2_valid & &tail ?
                io_op_bits_base_vs2_valid : ~(&tail) & _T_963) : _T_963;	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      wire [9:0] _T_1045 = io_op_bits_active_vfdiv ? (_T_132 ? io_op_bits_fn_union : _T_4 ? _T_1004 : _T_916) : _T_916;	// sequencer-master.scala:289:23
      wire [9:0] _T_1046 = io_op_bits_active_vfdiv ? (_T_133 ? io_op_bits_fn_union : _T_5 ? _T_1004 : _T_917) : _T_917;	// sequencer-master.scala:289:23
      wire [9:0] _T_1047 = io_op_bits_active_vfdiv ? (_T_134 ? io_op_bits_fn_union : _T_6 ? _T_1004 : _T_918) : _T_918;	// sequencer-master.scala:289:23
      wire [9:0] _T_1048 = io_op_bits_active_vfdiv ? (_T_135 ? io_op_bits_fn_union : _T_7 ? _T_1004 : _T_919) : _T_919;	// sequencer-master.scala:289:23
      wire [9:0] _T_1049 = io_op_bits_active_vfdiv ? (_T_136 ? io_op_bits_fn_union : _T_8 ? _T_1004 : _T_920) : _T_920;	// sequencer-master.scala:289:23
      wire [9:0] _T_1050 = io_op_bits_active_vfdiv ? (_T_137 ? io_op_bits_fn_union : _T_9 ? _T_1004 : _T_921) : _T_921;	// sequencer-master.scala:289:23
      wire [9:0] _T_1051 = io_op_bits_active_vfdiv ? (_T_138 ? io_op_bits_fn_union : _T_10 ? _T_1004 : _T_922) :
                _T_922;	// sequencer-master.scala:289:23
      wire [9:0] _T_1052 = io_op_bits_active_vfdiv ? (&_T_0 ? io_op_bits_fn_union : &tail ? _T_1004 : _T_923) : _T_923;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire [7:0] _T_1053 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_132 | _T_964 ?
                io_op_bits_base_vd_id : _T_876) : _T_964 ? io_op_bits_base_vd_id : _T_876;	// sequencer-master.scala:363:24
      wire _T_1054 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_132 ? io_op_bits_base_vd_valid :
                ~_T_132 & ~_T_4 & _T_965) : _T_965;	// sequencer-master.scala:276:28, :363:24
      wire _T_1055 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_132 | _T_966 ?
                io_op_bits_base_vd_scalar : _T_878) : _T_966 ? io_op_bits_base_vd_scalar : _T_878;	// sequencer-master.scala:363:24
      wire _T_1056 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_132 | _T_967 ?
                io_op_bits_base_vd_pred : _T_879) : _T_967 ? io_op_bits_base_vd_pred : _T_879;	// sequencer-master.scala:363:24
      wire [1:0] _T_1057 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_132 | _T_968 ?
                io_op_bits_base_vd_prec : _T_880) : _T_968 ? io_op_bits_base_vd_prec : _T_880;	// sequencer-master.scala:363:24
      wire [7:0] _T_1058 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_133 | _T_969 ?
                io_op_bits_base_vd_id : _T_881) : _T_969 ? io_op_bits_base_vd_id : _T_881;	// sequencer-master.scala:363:24
      wire _T_1059 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_133 ? io_op_bits_base_vd_valid :
                ~_T_133 & ~_T_5 & _T_970) : _T_970;	// sequencer-master.scala:276:28, :363:24
      wire _T_1060 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_133 | _T_971 ?
                io_op_bits_base_vd_scalar : _T_883) : _T_971 ? io_op_bits_base_vd_scalar : _T_883;	// sequencer-master.scala:363:24
      wire _T_1061 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_133 | _T_972 ?
                io_op_bits_base_vd_pred : _T_884) : _T_972 ? io_op_bits_base_vd_pred : _T_884;	// sequencer-master.scala:363:24
      wire [1:0] _T_1062 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_133 | _T_973 ?
                io_op_bits_base_vd_prec : _T_885) : _T_973 ? io_op_bits_base_vd_prec : _T_885;	// sequencer-master.scala:363:24
      wire [7:0] _T_1063 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_134 | _T_974 ?
                io_op_bits_base_vd_id : _T_886) : _T_974 ? io_op_bits_base_vd_id : _T_886;	// sequencer-master.scala:363:24
      wire _T_1064 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_134 ? io_op_bits_base_vd_valid :
                ~_T_134 & ~_T_6 & _T_975) : _T_975;	// sequencer-master.scala:276:28, :363:24
      wire _T_1065 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_134 | _T_976 ?
                io_op_bits_base_vd_scalar : _T_888) : _T_976 ? io_op_bits_base_vd_scalar : _T_888;	// sequencer-master.scala:363:24
      wire _T_1066 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_134 | _T_977 ?
                io_op_bits_base_vd_pred : _T_889) : _T_977 ? io_op_bits_base_vd_pred : _T_889;	// sequencer-master.scala:363:24
      wire [1:0] _T_1067 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_134 | _T_978 ?
                io_op_bits_base_vd_prec : _T_890) : _T_978 ? io_op_bits_base_vd_prec : _T_890;	// sequencer-master.scala:363:24
      wire [7:0] _T_1068 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_135 | _T_979 ?
                io_op_bits_base_vd_id : _T_891) : _T_979 ? io_op_bits_base_vd_id : _T_891;	// sequencer-master.scala:363:24
      wire _T_1069 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_135 ? io_op_bits_base_vd_valid :
                ~_T_135 & ~_T_7 & _T_980) : _T_980;	// sequencer-master.scala:276:28, :363:24
      wire _T_1070 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_135 | _T_981 ?
                io_op_bits_base_vd_scalar : _T_893) : _T_981 ? io_op_bits_base_vd_scalar : _T_893;	// sequencer-master.scala:363:24
      wire _T_1071 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_135 | _T_982 ?
                io_op_bits_base_vd_pred : _T_894) : _T_982 ? io_op_bits_base_vd_pred : _T_894;	// sequencer-master.scala:363:24
      wire [1:0] _T_1072 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_135 | _T_983 ?
                io_op_bits_base_vd_prec : _T_895) : _T_983 ? io_op_bits_base_vd_prec : _T_895;	// sequencer-master.scala:363:24
      wire [7:0] _T_1073 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_136 | _T_984 ?
                io_op_bits_base_vd_id : _T_896) : _T_984 ? io_op_bits_base_vd_id : _T_896;	// sequencer-master.scala:363:24
      wire _T_1074 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_136 ? io_op_bits_base_vd_valid :
                ~_T_136 & ~_T_8 & _T_985) : _T_985;	// sequencer-master.scala:276:28, :363:24
      wire _T_1075 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_136 | _T_986 ?
                io_op_bits_base_vd_scalar : _T_898) : _T_986 ? io_op_bits_base_vd_scalar : _T_898;	// sequencer-master.scala:363:24
      wire _T_1076 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_136 | _T_987 ?
                io_op_bits_base_vd_pred : _T_899) : _T_987 ? io_op_bits_base_vd_pred : _T_899;	// sequencer-master.scala:363:24
      wire [1:0] _T_1077 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_136 | _T_988 ?
                io_op_bits_base_vd_prec : _T_900) : _T_988 ? io_op_bits_base_vd_prec : _T_900;	// sequencer-master.scala:363:24
      wire [7:0] _T_1078 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_137 | _T_989 ?
                io_op_bits_base_vd_id : _T_901) : _T_989 ? io_op_bits_base_vd_id : _T_901;	// sequencer-master.scala:363:24
      wire _T_1079 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_137 ? io_op_bits_base_vd_valid :
                ~_T_137 & ~_T_9 & _T_990) : _T_990;	// sequencer-master.scala:276:28, :363:24
      wire _T_1080 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_137 | _T_991 ?
                io_op_bits_base_vd_scalar : _T_903) : _T_991 ? io_op_bits_base_vd_scalar : _T_903;	// sequencer-master.scala:363:24
      wire _T_1081 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_137 | _T_992 ?
                io_op_bits_base_vd_pred : _T_904) : _T_992 ? io_op_bits_base_vd_pred : _T_904;	// sequencer-master.scala:363:24
      wire [1:0] _T_1082 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_137 | _T_993 ?
                io_op_bits_base_vd_prec : _T_905) : _T_993 ? io_op_bits_base_vd_prec : _T_905;	// sequencer-master.scala:363:24
      wire [7:0] _T_1083 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_138 | _T_994 ?
                io_op_bits_base_vd_id : _T_906) : _T_994 ? io_op_bits_base_vd_id : _T_906;	// sequencer-master.scala:363:24
      wire _T_1084 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & _T_138 ? io_op_bits_base_vd_valid :
                ~_T_138 & ~_T_10 & _T_995) : _T_995;	// sequencer-master.scala:276:28, :363:24
      wire _T_1085 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_138 | _T_996 ?
                io_op_bits_base_vd_scalar : _T_908) : _T_996 ? io_op_bits_base_vd_scalar : _T_908;	// sequencer-master.scala:363:24
      wire _T_1086 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_138 | _T_997 ?
                io_op_bits_base_vd_pred : _T_909) : _T_997 ? io_op_bits_base_vd_pred : _T_909;	// sequencer-master.scala:363:24
      wire [1:0] _T_1087 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (_T_138 | _T_998 ?
                io_op_bits_base_vd_prec : _T_910) : _T_998 ? io_op_bits_base_vd_prec : _T_910;	// sequencer-master.scala:363:24
      wire [7:0] _T_1088 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_999 ?
                io_op_bits_base_vd_id : _T_911) : _T_999 ? io_op_bits_base_vd_id : _T_911;	// sequencer-master.scala:267:35, :363:24
      wire _T_1089 = io_op_bits_active_vfdiv ? (io_op_bits_base_vd_valid & &_T_0 ? io_op_bits_base_vd_valid :
                ~(&_T_0) & ~(&tail) & _T_1000) : _T_1000;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_1090 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_1001 ?
                io_op_bits_base_vd_scalar : _T_913) : _T_1001 ? io_op_bits_base_vd_scalar : _T_913;	// sequencer-master.scala:267:35, :363:24
      wire _T_1091 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_1002 ?
                io_op_bits_base_vd_pred : _T_914) : _T_1002 ? io_op_bits_base_vd_pred : _T_914;	// sequencer-master.scala:267:35, :363:24
      wire [1:0] _T_1092 = io_op_bits_active_vfdiv & io_op_bits_base_vd_valid ? (&_T_0 | _T_1003 ?
                io_op_bits_base_vd_prec : _T_915) : _T_1003 ? io_op_bits_base_vd_prec : _T_915;	// sequencer-master.scala:267:35, :363:24
      wire _T_1093 = io_op_bits_active_vfcmp & _T_4;	// sequencer-master.scala:289:23
      wire _T_1094 = io_op_bits_active_vfcmp & _T_5;	// sequencer-master.scala:289:23
      wire _T_1095 = io_op_bits_active_vfcmp & _T_6;	// sequencer-master.scala:289:23
      wire _T_1096 = io_op_bits_active_vfcmp & _T_7;	// sequencer-master.scala:289:23
      wire _T_1097 = io_op_bits_active_vfcmp & _T_8;	// sequencer-master.scala:289:23
      wire _T_1098 = io_op_bits_active_vfcmp & _T_9;	// sequencer-master.scala:289:23
      wire _T_1099 = io_op_bits_active_vfcmp & _T_10;	// sequencer-master.scala:289:23
      wire _T_1100 = io_op_bits_active_vfcmp & &tail;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire [3:0] _T_1101 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_4 | _T_1005 ?
                io_op_bits_base_vp_id : _T_924) : _T_1005 ? io_op_bits_base_vp_id : _T_924;	// sequencer-master.scala:321:24
      wire _T_1102 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_1029) : _T_1029;	// sequencer-master.scala:272:28, :321:24
      wire _T_1103 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_4 | _T_1006 ?
                io_op_bits_base_vp_scalar : _T_926) : _T_1006 ? io_op_bits_base_vp_scalar : _T_926;	// sequencer-master.scala:321:24
      wire _T_1104 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_4 | _T_1007 ?
                io_op_bits_base_vp_pred : _T_927) : _T_1007 ? io_op_bits_base_vp_pred : _T_927;	// sequencer-master.scala:321:24
      wire [3:0] _T_1105 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_5 | _T_1008 ?
                io_op_bits_base_vp_id : _T_928) : _T_1008 ? io_op_bits_base_vp_id : _T_928;	// sequencer-master.scala:321:24
      wire _T_1106 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_1030) : _T_1030;	// sequencer-master.scala:272:28, :321:24
      wire _T_1107 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_5 | _T_1009 ?
                io_op_bits_base_vp_scalar : _T_930) : _T_1009 ? io_op_bits_base_vp_scalar : _T_930;	// sequencer-master.scala:321:24
      wire _T_1108 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_5 | _T_1010 ?
                io_op_bits_base_vp_pred : _T_931) : _T_1010 ? io_op_bits_base_vp_pred : _T_931;	// sequencer-master.scala:321:24
      wire [3:0] _T_1109 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_6 | _T_1011 ?
                io_op_bits_base_vp_id : _T_932) : _T_1011 ? io_op_bits_base_vp_id : _T_932;	// sequencer-master.scala:321:24
      wire _T_1110 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_1031) : _T_1031;	// sequencer-master.scala:272:28, :321:24
      wire _T_1111 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_6 | _T_1012 ?
                io_op_bits_base_vp_scalar : _T_934) : _T_1012 ? io_op_bits_base_vp_scalar : _T_934;	// sequencer-master.scala:321:24
      wire _T_1112 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_6 | _T_1013 ?
                io_op_bits_base_vp_pred : _T_935) : _T_1013 ? io_op_bits_base_vp_pred : _T_935;	// sequencer-master.scala:321:24
      wire [3:0] _T_1113 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_7 | _T_1014 ?
                io_op_bits_base_vp_id : _T_936) : _T_1014 ? io_op_bits_base_vp_id : _T_936;	// sequencer-master.scala:321:24
      wire _T_1114 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_1032) : _T_1032;	// sequencer-master.scala:272:28, :321:24
      wire _T_1115 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_7 | _T_1015 ?
                io_op_bits_base_vp_scalar : _T_938) : _T_1015 ? io_op_bits_base_vp_scalar : _T_938;	// sequencer-master.scala:321:24
      wire _T_1116 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_7 | _T_1016 ?
                io_op_bits_base_vp_pred : _T_939) : _T_1016 ? io_op_bits_base_vp_pred : _T_939;	// sequencer-master.scala:321:24
      wire [3:0] _T_1117 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_8 | _T_1017 ?
                io_op_bits_base_vp_id : _T_940) : _T_1017 ? io_op_bits_base_vp_id : _T_940;	// sequencer-master.scala:321:24
      wire _T_1118 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_1033) : _T_1033;	// sequencer-master.scala:272:28, :321:24
      wire _T_1119 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_8 | _T_1018 ?
                io_op_bits_base_vp_scalar : _T_942) : _T_1018 ? io_op_bits_base_vp_scalar : _T_942;	// sequencer-master.scala:321:24
      wire _T_1120 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_8 | _T_1019 ?
                io_op_bits_base_vp_pred : _T_943) : _T_1019 ? io_op_bits_base_vp_pred : _T_943;	// sequencer-master.scala:321:24
      wire [3:0] _T_1121 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_9 | _T_1020 ?
                io_op_bits_base_vp_id : _T_944) : _T_1020 ? io_op_bits_base_vp_id : _T_944;	// sequencer-master.scala:321:24
      wire _T_1122 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_1034) : _T_1034;	// sequencer-master.scala:272:28, :321:24
      wire _T_1123 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_9 | _T_1021 ?
                io_op_bits_base_vp_scalar : _T_946) : _T_1021 ? io_op_bits_base_vp_scalar : _T_946;	// sequencer-master.scala:321:24
      wire _T_1124 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_9 | _T_1022 ?
                io_op_bits_base_vp_pred : _T_947) : _T_1022 ? io_op_bits_base_vp_pred : _T_947;	// sequencer-master.scala:321:24
      wire [3:0] _T_1125 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_10 | _T_1023 ?
                io_op_bits_base_vp_id : _T_948) : _T_1023 ? io_op_bits_base_vp_id : _T_948;	// sequencer-master.scala:321:24
      wire _T_1126 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_1035) : _T_1035;	// sequencer-master.scala:272:28, :321:24
      wire _T_1127 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_10 | _T_1024 ?
                io_op_bits_base_vp_scalar : _T_950) : _T_1024 ? io_op_bits_base_vp_scalar : _T_950;	// sequencer-master.scala:321:24
      wire _T_1128 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (_T_10 | _T_1025 ?
                io_op_bits_base_vp_pred : _T_951) : _T_1025 ? io_op_bits_base_vp_pred : _T_951;	// sequencer-master.scala:321:24
      wire [3:0] _T_1129 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (&tail | _T_1026 ?
                io_op_bits_base_vp_id : _T_952) : _T_1026 ? io_op_bits_base_vp_id : _T_952;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1130 = io_op_bits_active_vfcmp ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_1036) : _T_1036;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1131 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (&tail | _T_1027 ?
                io_op_bits_base_vp_scalar : _T_954) : _T_1027 ? io_op_bits_base_vp_scalar : _T_954;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1132 = io_op_bits_active_vfcmp & io_op_bits_base_vp_valid ? (&tail | _T_1028 ?
                io_op_bits_base_vp_pred : _T_955) : _T_1028 ? io_op_bits_base_vp_pred : _T_955;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1133 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_1134 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & _T_1054) : _T_1054;	// sequencer-master.scala:276:28, :363:24
      wire _T_1135 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_1136 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_1137 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_4;	// sequencer-master.scala:363:24
      wire _T_1138 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_1139 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & _T_1059) : _T_1059;	// sequencer-master.scala:276:28, :363:24
      wire _T_1140 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_1141 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_1142 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_5;	// sequencer-master.scala:363:24
      wire _T_1143 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_1144 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & _T_1064) : _T_1064;	// sequencer-master.scala:276:28, :363:24
      wire _T_1145 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_1146 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_1147 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_6;	// sequencer-master.scala:363:24
      wire _T_1148 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_1149 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & _T_1069) : _T_1069;	// sequencer-master.scala:276:28, :363:24
      wire _T_1150 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_1151 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_1152 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_7;	// sequencer-master.scala:363:24
      wire _T_1153 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_1154 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & _T_1074) : _T_1074;	// sequencer-master.scala:276:28, :363:24
      wire _T_1155 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_1156 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_1157 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_8;	// sequencer-master.scala:363:24
      wire _T_1158 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_1159 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & _T_1079) : _T_1079;	// sequencer-master.scala:276:28, :363:24
      wire _T_1160 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_1161 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_1162 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_9;	// sequencer-master.scala:363:24
      wire _T_1163 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_1164 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & _T_1084) : _T_1084;	// sequencer-master.scala:276:28, :363:24
      wire _T_1165 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_1166 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_1167 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & _T_10;	// sequencer-master.scala:363:24
      wire _T_1168 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1169 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & _T_1089) : _T_1089;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_1170 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1171 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1172 = io_op_bits_active_vfcmp & io_op_bits_base_vd_valid & &tail;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1173 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1174 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_1102) : _T_1102;	// sequencer-master.scala:272:28, :321:24
      wire _T_1175 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1176 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1177 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1178 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_1106) : _T_1106;	// sequencer-master.scala:272:28, :321:24
      wire _T_1179 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1180 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1181 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1182 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_1110) : _T_1110;	// sequencer-master.scala:272:28, :321:24
      wire _T_1183 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1184 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1185 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1186 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_1114) : _T_1114;	// sequencer-master.scala:272:28, :321:24
      wire _T_1187 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1188 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1189 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1190 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_1118) : _T_1118;	// sequencer-master.scala:272:28, :321:24
      wire _T_1191 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1192 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1193 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1194 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_1122) : _T_1122;	// sequencer-master.scala:272:28, :321:24
      wire _T_1195 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1196 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1197 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1198 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_1126) : _T_1126;	// sequencer-master.scala:272:28, :321:24
      wire _T_1199 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1200 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1201 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1202 = io_op_bits_active_vfconv ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_1130) : _T_1130;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1203 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1204 = io_op_bits_active_vfconv & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire [7:0] _T_1205 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_4 | _T_1133 ?
                io_op_bits_base_vd_id : _T_1053) : _T_1133 ? io_op_bits_base_vd_id : _T_1053;	// sequencer-master.scala:363:24
      wire _T_1206 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_4 | _T_1135 ?
                io_op_bits_base_vd_scalar : _T_1055) : _T_1135 ? io_op_bits_base_vd_scalar : _T_1055;	// sequencer-master.scala:363:24
      wire _T_1207 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_4 | _T_1136 ?
                io_op_bits_base_vd_pred : _T_1056) : _T_1136 ? io_op_bits_base_vd_pred : _T_1056;	// sequencer-master.scala:363:24
      wire [1:0] _T_1208 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_4 | _T_1137 ?
                io_op_bits_base_vd_prec : _T_1057) : _T_1137 ? io_op_bits_base_vd_prec : _T_1057;	// sequencer-master.scala:363:24
      wire [7:0] _T_1209 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_5 | _T_1138 ?
                io_op_bits_base_vd_id : _T_1058) : _T_1138 ? io_op_bits_base_vd_id : _T_1058;	// sequencer-master.scala:363:24
      wire _T_1210 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_5 | _T_1140 ?
                io_op_bits_base_vd_scalar : _T_1060) : _T_1140 ? io_op_bits_base_vd_scalar : _T_1060;	// sequencer-master.scala:363:24
      wire _T_1211 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_5 | _T_1141 ?
                io_op_bits_base_vd_pred : _T_1061) : _T_1141 ? io_op_bits_base_vd_pred : _T_1061;	// sequencer-master.scala:363:24
      wire [1:0] _T_1212 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_5 | _T_1142 ?
                io_op_bits_base_vd_prec : _T_1062) : _T_1142 ? io_op_bits_base_vd_prec : _T_1062;	// sequencer-master.scala:363:24
      wire [7:0] _T_1213 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_6 | _T_1143 ?
                io_op_bits_base_vd_id : _T_1063) : _T_1143 ? io_op_bits_base_vd_id : _T_1063;	// sequencer-master.scala:363:24
      wire _T_1214 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_6 | _T_1145 ?
                io_op_bits_base_vd_scalar : _T_1065) : _T_1145 ? io_op_bits_base_vd_scalar : _T_1065;	// sequencer-master.scala:363:24
      wire _T_1215 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_6 | _T_1146 ?
                io_op_bits_base_vd_pred : _T_1066) : _T_1146 ? io_op_bits_base_vd_pred : _T_1066;	// sequencer-master.scala:363:24
      wire [1:0] _T_1216 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_6 | _T_1147 ?
                io_op_bits_base_vd_prec : _T_1067) : _T_1147 ? io_op_bits_base_vd_prec : _T_1067;	// sequencer-master.scala:363:24
      wire [7:0] _T_1217 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_7 | _T_1148 ?
                io_op_bits_base_vd_id : _T_1068) : _T_1148 ? io_op_bits_base_vd_id : _T_1068;	// sequencer-master.scala:363:24
      wire _T_1218 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_7 | _T_1150 ?
                io_op_bits_base_vd_scalar : _T_1070) : _T_1150 ? io_op_bits_base_vd_scalar : _T_1070;	// sequencer-master.scala:363:24
      wire _T_1219 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_7 | _T_1151 ?
                io_op_bits_base_vd_pred : _T_1071) : _T_1151 ? io_op_bits_base_vd_pred : _T_1071;	// sequencer-master.scala:363:24
      wire [1:0] _T_1220 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_7 | _T_1152 ?
                io_op_bits_base_vd_prec : _T_1072) : _T_1152 ? io_op_bits_base_vd_prec : _T_1072;	// sequencer-master.scala:363:24
      wire [7:0] _T_1221 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_8 | _T_1153 ?
                io_op_bits_base_vd_id : _T_1073) : _T_1153 ? io_op_bits_base_vd_id : _T_1073;	// sequencer-master.scala:363:24
      wire _T_1222 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_8 | _T_1155 ?
                io_op_bits_base_vd_scalar : _T_1075) : _T_1155 ? io_op_bits_base_vd_scalar : _T_1075;	// sequencer-master.scala:363:24
      wire _T_1223 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_8 | _T_1156 ?
                io_op_bits_base_vd_pred : _T_1076) : _T_1156 ? io_op_bits_base_vd_pred : _T_1076;	// sequencer-master.scala:363:24
      wire [1:0] _T_1224 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_8 | _T_1157 ?
                io_op_bits_base_vd_prec : _T_1077) : _T_1157 ? io_op_bits_base_vd_prec : _T_1077;	// sequencer-master.scala:363:24
      wire [7:0] _T_1225 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_9 | _T_1158 ?
                io_op_bits_base_vd_id : _T_1078) : _T_1158 ? io_op_bits_base_vd_id : _T_1078;	// sequencer-master.scala:363:24
      wire _T_1226 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_9 | _T_1160 ?
                io_op_bits_base_vd_scalar : _T_1080) : _T_1160 ? io_op_bits_base_vd_scalar : _T_1080;	// sequencer-master.scala:363:24
      wire _T_1227 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_9 | _T_1161 ?
                io_op_bits_base_vd_pred : _T_1081) : _T_1161 ? io_op_bits_base_vd_pred : _T_1081;	// sequencer-master.scala:363:24
      wire [1:0] _T_1228 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_9 | _T_1162 ?
                io_op_bits_base_vd_prec : _T_1082) : _T_1162 ? io_op_bits_base_vd_prec : _T_1082;	// sequencer-master.scala:363:24
      wire [7:0] _T_1229 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_10 | _T_1163 ?
                io_op_bits_base_vd_id : _T_1083) : _T_1163 ? io_op_bits_base_vd_id : _T_1083;	// sequencer-master.scala:363:24
      wire _T_1230 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_10 | _T_1165 ?
                io_op_bits_base_vd_scalar : _T_1085) : _T_1165 ? io_op_bits_base_vd_scalar : _T_1085;	// sequencer-master.scala:363:24
      wire _T_1231 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_10 | _T_1166 ?
                io_op_bits_base_vd_pred : _T_1086) : _T_1166 ? io_op_bits_base_vd_pred : _T_1086;	// sequencer-master.scala:363:24
      wire [1:0] _T_1232 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (_T_10 | _T_1167 ?
                io_op_bits_base_vd_prec : _T_1087) : _T_1167 ? io_op_bits_base_vd_prec : _T_1087;	// sequencer-master.scala:363:24
      wire [7:0] _T_1233 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (&tail | _T_1168 ?
                io_op_bits_base_vd_id : _T_1088) : _T_1168 ? io_op_bits_base_vd_id : _T_1088;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1234 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (&tail | _T_1170 ?
                io_op_bits_base_vd_scalar : _T_1090) : _T_1170 ? io_op_bits_base_vd_scalar : _T_1090;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire _T_1235 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (&tail | _T_1171 ?
                io_op_bits_base_vd_pred : _T_1091) : _T_1171 ? io_op_bits_base_vd_pred : _T_1091;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire [1:0] _T_1236 = io_op_bits_active_vfconv & io_op_bits_base_vd_valid ? (&tail | _T_1172 ?
                io_op_bits_base_vd_prec : _T_1092) : _T_1172 ? io_op_bits_base_vd_prec : _T_1092;	// sequencer-master.scala:267:35, :363:24, util.scala:94:11
      wire [9:0] _T_1237 = {8'h0, io_op_bits_active_vidiv | io_op_bits_active_vfdiv & ~(io_op_bits_fn_union[0]),
                _T_826};	// sequencer-master.scala:289:23, :300:{28,46}, :411:70, types-vxu.scala:54:51, :96:47
      wire [3:0] _T_1238 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_4 | _T_1173 ?
                io_op_bits_base_vp_id : _T_1101) : _T_1173 ? io_op_bits_base_vp_id : _T_1101;	// sequencer-master.scala:321:24
      wire _T_1239 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_1174) : _T_1174;	// sequencer-master.scala:272:28, :321:24
      wire _T_1240 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_4 | _T_1175 ?
                io_op_bits_base_vp_scalar : _T_1103) : _T_1175 ? io_op_bits_base_vp_scalar : _T_1103;	// sequencer-master.scala:321:24
      wire _T_1241 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_4 | _T_1176 ?
                io_op_bits_base_vp_pred : _T_1104) : _T_1176 ? io_op_bits_base_vp_pred : _T_1104;	// sequencer-master.scala:321:24
      wire [3:0] _T_1242 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_5 | _T_1177 ?
                io_op_bits_base_vp_id : _T_1105) : _T_1177 ? io_op_bits_base_vp_id : _T_1105;	// sequencer-master.scala:321:24
      wire _T_1243 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_1178) : _T_1178;	// sequencer-master.scala:272:28, :321:24
      wire _T_1244 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_5 | _T_1179 ?
                io_op_bits_base_vp_scalar : _T_1107) : _T_1179 ? io_op_bits_base_vp_scalar : _T_1107;	// sequencer-master.scala:321:24
      wire _T_1245 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_5 | _T_1180 ?
                io_op_bits_base_vp_pred : _T_1108) : _T_1180 ? io_op_bits_base_vp_pred : _T_1108;	// sequencer-master.scala:321:24
      wire [3:0] _T_1246 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_6 | _T_1181 ?
                io_op_bits_base_vp_id : _T_1109) : _T_1181 ? io_op_bits_base_vp_id : _T_1109;	// sequencer-master.scala:321:24
      wire _T_1247 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_1182) : _T_1182;	// sequencer-master.scala:272:28, :321:24
      wire _T_1248 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_6 | _T_1183 ?
                io_op_bits_base_vp_scalar : _T_1111) : _T_1183 ? io_op_bits_base_vp_scalar : _T_1111;	// sequencer-master.scala:321:24
      wire _T_1249 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_6 | _T_1184 ?
                io_op_bits_base_vp_pred : _T_1112) : _T_1184 ? io_op_bits_base_vp_pred : _T_1112;	// sequencer-master.scala:321:24
      wire [3:0] _T_1250 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_7 | _T_1185 ?
                io_op_bits_base_vp_id : _T_1113) : _T_1185 ? io_op_bits_base_vp_id : _T_1113;	// sequencer-master.scala:321:24
      wire _T_1251 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_1186) : _T_1186;	// sequencer-master.scala:272:28, :321:24
      wire _T_1252 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_7 | _T_1187 ?
                io_op_bits_base_vp_scalar : _T_1115) : _T_1187 ? io_op_bits_base_vp_scalar : _T_1115;	// sequencer-master.scala:321:24
      wire _T_1253 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_7 | _T_1188 ?
                io_op_bits_base_vp_pred : _T_1116) : _T_1188 ? io_op_bits_base_vp_pred : _T_1116;	// sequencer-master.scala:321:24
      wire [3:0] _T_1254 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_8 | _T_1189 ?
                io_op_bits_base_vp_id : _T_1117) : _T_1189 ? io_op_bits_base_vp_id : _T_1117;	// sequencer-master.scala:321:24
      wire _T_1255 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_1190) : _T_1190;	// sequencer-master.scala:272:28, :321:24
      wire _T_1256 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_8 | _T_1191 ?
                io_op_bits_base_vp_scalar : _T_1119) : _T_1191 ? io_op_bits_base_vp_scalar : _T_1119;	// sequencer-master.scala:321:24
      wire _T_1257 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_8 | _T_1192 ?
                io_op_bits_base_vp_pred : _T_1120) : _T_1192 ? io_op_bits_base_vp_pred : _T_1120;	// sequencer-master.scala:321:24
      wire [3:0] _T_1258 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_9 | _T_1193 ?
                io_op_bits_base_vp_id : _T_1121) : _T_1193 ? io_op_bits_base_vp_id : _T_1121;	// sequencer-master.scala:321:24
      wire _T_1259 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_1194) : _T_1194;	// sequencer-master.scala:272:28, :321:24
      wire _T_1260 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_9 | _T_1195 ?
                io_op_bits_base_vp_scalar : _T_1123) : _T_1195 ? io_op_bits_base_vp_scalar : _T_1123;	// sequencer-master.scala:321:24
      wire _T_1261 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_9 | _T_1196 ?
                io_op_bits_base_vp_pred : _T_1124) : _T_1196 ? io_op_bits_base_vp_pred : _T_1124;	// sequencer-master.scala:321:24
      wire [3:0] _T_1262 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_10 | _T_1197 ?
                io_op_bits_base_vp_id : _T_1125) : _T_1197 ? io_op_bits_base_vp_id : _T_1125;	// sequencer-master.scala:321:24
      wire _T_1263 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_1198) : _T_1198;	// sequencer-master.scala:272:28, :321:24
      wire _T_1264 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_10 | _T_1199 ?
                io_op_bits_base_vp_scalar : _T_1127) : _T_1199 ? io_op_bits_base_vp_scalar : _T_1127;	// sequencer-master.scala:321:24
      wire _T_1265 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (_T_10 | _T_1200 ?
                io_op_bits_base_vp_pred : _T_1128) : _T_1200 ? io_op_bits_base_vp_pred : _T_1128;	// sequencer-master.scala:321:24
      wire [3:0] _T_1266 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (&tail | _T_1201 ?
                io_op_bits_base_vp_id : _T_1129) : _T_1201 ? io_op_bits_base_vp_id : _T_1129;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1267 = io_op_bits_active_vrpred ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_1202) : _T_1202;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1268 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (&tail | _T_1203 ?
                io_op_bits_base_vp_scalar : _T_1131) : _T_1203 ? io_op_bits_base_vp_scalar : _T_1131;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1269 = io_op_bits_active_vrpred & io_op_bits_base_vp_valid ? (&tail | _T_1204 ?
                io_op_bits_base_vp_pred : _T_1132) : _T_1204 ? io_op_bits_base_vp_pred : _T_1132;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1270 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_4 ? io_op_bits_base_vd_valid :
                ~_T_4 & _T_1134) : _T_1134);	// sequencer-master.scala:276:28, :363:24
      wire _T_1271 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_5 ? io_op_bits_base_vd_valid :
                ~_T_5 & _T_1139) : _T_1139);	// sequencer-master.scala:276:28, :363:24
      wire _T_1272 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_6 ? io_op_bits_base_vd_valid :
                ~_T_6 & _T_1144) : _T_1144);	// sequencer-master.scala:276:28, :363:24
      wire _T_1273 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_7 ? io_op_bits_base_vd_valid :
                ~_T_7 & _T_1149) : _T_1149);	// sequencer-master.scala:276:28, :363:24
      wire _T_1274 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_8 ? io_op_bits_base_vd_valid :
                ~_T_8 & _T_1154) : _T_1154);	// sequencer-master.scala:276:28, :363:24
      wire _T_1275 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_9 ? io_op_bits_base_vd_valid :
                ~_T_9 & _T_1159) : _T_1159);	// sequencer-master.scala:276:28, :363:24
      wire _T_1276 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & _T_10 ? io_op_bits_base_vd_valid :
                ~_T_10 & _T_1164) : _T_1164);	// sequencer-master.scala:276:28, :363:24
      wire _T_1277 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? (io_op_bits_base_vd_valid & &tail ? io_op_bits_base_vd_valid :
                ~(&tail) & _T_1169) : _T_1169);	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire [9:0] _T_1278 = {8'h0, io_op_bits_active_vidiv | io_op_bits_active_vfdiv & ~(io_op_bits_fn_union[0]),
                _T_826};	// sequencer-master.scala:289:23, :300:{28,46}, :411:70, types-vxu.scala:54:51, :96:47
      wire [9:0] _T_1279 = io_op_bits_active_vrfirst & _T_4 ? _T_1278 : io_op_bits_active_vrpred & _T_4 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_4 | _T_1093 ? io_op_bits_fn_union : _T_1045) : _T_1093 ?
                io_op_bits_fn_union : _T_1045;	// sequencer-master.scala:289:23
      wire [9:0] _T_1280 = io_op_bits_active_vrfirst & _T_5 ? _T_1278 : io_op_bits_active_vrpred & _T_5 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_5 | _T_1094 ? io_op_bits_fn_union : _T_1046) : _T_1094 ?
                io_op_bits_fn_union : _T_1046;	// sequencer-master.scala:289:23
      wire [9:0] _T_1281 = io_op_bits_active_vrfirst & _T_6 ? _T_1278 : io_op_bits_active_vrpred & _T_6 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_6 | _T_1095 ? io_op_bits_fn_union : _T_1047) : _T_1095 ?
                io_op_bits_fn_union : _T_1047;	// sequencer-master.scala:289:23
      wire [9:0] _T_1282 = io_op_bits_active_vrfirst & _T_7 ? _T_1278 : io_op_bits_active_vrpred & _T_7 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_7 | _T_1096 ? io_op_bits_fn_union : _T_1048) : _T_1096 ?
                io_op_bits_fn_union : _T_1048;	// sequencer-master.scala:289:23
      wire [9:0] _T_1283 = io_op_bits_active_vrfirst & _T_8 ? _T_1278 : io_op_bits_active_vrpred & _T_8 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_8 | _T_1097 ? io_op_bits_fn_union : _T_1049) : _T_1097 ?
                io_op_bits_fn_union : _T_1049;	// sequencer-master.scala:289:23
      wire [9:0] _T_1284 = io_op_bits_active_vrfirst & _T_9 ? _T_1278 : io_op_bits_active_vrpred & _T_9 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_9 | _T_1098 ? io_op_bits_fn_union : _T_1050) : _T_1098 ?
                io_op_bits_fn_union : _T_1050;	// sequencer-master.scala:289:23
      wire [9:0] _T_1285 = io_op_bits_active_vrfirst & _T_10 ? _T_1278 : io_op_bits_active_vrpred & _T_10 ? _T_1237 :
                io_op_bits_active_vfconv ? (_T_10 | _T_1099 ? io_op_bits_fn_union : _T_1051) : _T_1099 ?
                io_op_bits_fn_union : _T_1051;	// sequencer-master.scala:289:23
      wire [9:0] _T_1286 = io_op_bits_active_vrfirst & &tail ? _T_1278 : io_op_bits_active_vrpred & &tail ? _T_1237 :
                io_op_bits_active_vfconv ? (&tail | _T_1100 ? io_op_bits_fn_union : _T_1052) : _T_1100 ?
                io_op_bits_fn_union : _T_1052;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire _T_1287 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire [3:0] _T_1288 = _T_1287 ? io_op_bits_base_vp_id : _T_1238;	// sequencer-master.scala:321:24
      wire _T_1289 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid :
                ~_T_4 & _T_1239) : _T_1239;	// sequencer-master.scala:272:28, :321:24
      wire _T_1290 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1291 = _T_1290 ? io_op_bits_base_vp_scalar : _T_1240;	// sequencer-master.scala:321:24
      wire _T_1292 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1293 = _T_1292 ? io_op_bits_base_vp_pred : _T_1241;	// sequencer-master.scala:321:24
      wire _T_1294 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire [3:0] _T_1295 = _T_1294 ? io_op_bits_base_vp_id : _T_1242;	// sequencer-master.scala:321:24
      wire _T_1296 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid :
                ~_T_5 & _T_1243) : _T_1243;	// sequencer-master.scala:272:28, :321:24
      wire _T_1297 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1298 = _T_1297 ? io_op_bits_base_vp_scalar : _T_1244;	// sequencer-master.scala:321:24
      wire _T_1299 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1300 = _T_1299 ? io_op_bits_base_vp_pred : _T_1245;	// sequencer-master.scala:321:24
      wire _T_1301 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire [3:0] _T_1302 = _T_1301 ? io_op_bits_base_vp_id : _T_1246;	// sequencer-master.scala:321:24
      wire _T_1303 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid :
                ~_T_6 & _T_1247) : _T_1247;	// sequencer-master.scala:272:28, :321:24
      wire _T_1304 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1305 = _T_1304 ? io_op_bits_base_vp_scalar : _T_1248;	// sequencer-master.scala:321:24
      wire _T_1306 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1307 = _T_1306 ? io_op_bits_base_vp_pred : _T_1249;	// sequencer-master.scala:321:24
      wire _T_1308 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire [3:0] _T_1309 = _T_1308 ? io_op_bits_base_vp_id : _T_1250;	// sequencer-master.scala:321:24
      wire _T_1310 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid :
                ~_T_7 & _T_1251) : _T_1251;	// sequencer-master.scala:272:28, :321:24
      wire _T_1311 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1312 = _T_1311 ? io_op_bits_base_vp_scalar : _T_1252;	// sequencer-master.scala:321:24
      wire _T_1313 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1314 = _T_1313 ? io_op_bits_base_vp_pred : _T_1253;	// sequencer-master.scala:321:24
      wire _T_1315 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire [3:0] _T_1316 = _T_1315 ? io_op_bits_base_vp_id : _T_1254;	// sequencer-master.scala:321:24
      wire _T_1317 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid :
                ~_T_8 & _T_1255) : _T_1255;	// sequencer-master.scala:272:28, :321:24
      wire _T_1318 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1319 = _T_1318 ? io_op_bits_base_vp_scalar : _T_1256;	// sequencer-master.scala:321:24
      wire _T_1320 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1321 = _T_1320 ? io_op_bits_base_vp_pred : _T_1257;	// sequencer-master.scala:321:24
      wire _T_1322 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire [3:0] _T_1323 = _T_1322 ? io_op_bits_base_vp_id : _T_1258;	// sequencer-master.scala:321:24
      wire _T_1324 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid :
                ~_T_9 & _T_1259) : _T_1259;	// sequencer-master.scala:272:28, :321:24
      wire _T_1325 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1326 = _T_1325 ? io_op_bits_base_vp_scalar : _T_1260;	// sequencer-master.scala:321:24
      wire _T_1327 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1328 = _T_1327 ? io_op_bits_base_vp_pred : _T_1261;	// sequencer-master.scala:321:24
      wire _T_1329 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire [3:0] _T_1330 = _T_1329 ? io_op_bits_base_vp_id : _T_1262;	// sequencer-master.scala:321:24
      wire _T_1331 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid :
                ~_T_10 & _T_1263) : _T_1263;	// sequencer-master.scala:272:28, :321:24
      wire _T_1332 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1333 = _T_1332 ? io_op_bits_base_vp_scalar : _T_1264;	// sequencer-master.scala:321:24
      wire _T_1334 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1335 = _T_1334 ? io_op_bits_base_vp_pred : _T_1265;	// sequencer-master.scala:321:24
      wire _T_1336 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire [3:0] _T_1337 = _T_1336 ? io_op_bits_base_vp_id : _T_1266;	// sequencer-master.scala:321:24
      wire _T_1338 = io_op_bits_active_vrfirst ? (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_1267) : _T_1267;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1339 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1340 = _T_1339 ? io_op_bits_base_vp_scalar : _T_1268;	// sequencer-master.scala:321:24
      wire _T_1341 = io_op_bits_active_vrfirst & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1342 = _T_1341 ? io_op_bits_base_vp_pred : _T_1269;	// sequencer-master.scala:321:24
      wire [3:0] _T_1343 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1287 ? io_op_bits_base_vp_id : _T_1238) : _T_1288) :
                _T_1288;	// sequencer-master.scala:321:24
      wire _T_1344 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1290 ? io_op_bits_base_vp_scalar : _T_1240) :
                _T_1291) : _T_1291;	// sequencer-master.scala:321:24
      wire _T_1345 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1292 ? io_op_bits_base_vp_pred : _T_1241) : _T_1293)
                : _T_1293;	// sequencer-master.scala:321:24
      wire [3:0] _T_1346 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1294 ? io_op_bits_base_vp_id : _T_1242) : _T_1295) :
                _T_1295;	// sequencer-master.scala:321:24
      wire _T_1347 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1297 ? io_op_bits_base_vp_scalar : _T_1244) :
                _T_1298) : _T_1298;	// sequencer-master.scala:321:24
      wire _T_1348 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1299 ? io_op_bits_base_vp_pred : _T_1245) : _T_1300)
                : _T_1300;	// sequencer-master.scala:321:24
      wire [3:0] _T_1349 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1301 ? io_op_bits_base_vp_id : _T_1246) : _T_1302) :
                _T_1302;	// sequencer-master.scala:321:24
      wire _T_1350 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1304 ? io_op_bits_base_vp_scalar : _T_1248) :
                _T_1305) : _T_1305;	// sequencer-master.scala:321:24
      wire _T_1351 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1306 ? io_op_bits_base_vp_pred : _T_1249) : _T_1307)
                : _T_1307;	// sequencer-master.scala:321:24
      wire [3:0] _T_1352 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1308 ? io_op_bits_base_vp_id : _T_1250) : _T_1309) :
                _T_1309;	// sequencer-master.scala:321:24
      wire _T_1353 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1311 ? io_op_bits_base_vp_scalar : _T_1252) :
                _T_1312) : _T_1312;	// sequencer-master.scala:321:24
      wire _T_1354 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1313 ? io_op_bits_base_vp_pred : _T_1253) : _T_1314)
                : _T_1314;	// sequencer-master.scala:321:24
      wire [3:0] _T_1355 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1315 ? io_op_bits_base_vp_id : _T_1254) : _T_1316) :
                _T_1316;	// sequencer-master.scala:321:24
      wire _T_1356 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1318 ? io_op_bits_base_vp_scalar : _T_1256) :
                _T_1319) : _T_1319;	// sequencer-master.scala:321:24
      wire _T_1357 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1320 ? io_op_bits_base_vp_pred : _T_1257) : _T_1321)
                : _T_1321;	// sequencer-master.scala:321:24
      wire [3:0] _T_1358 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1322 ? io_op_bits_base_vp_id : _T_1258) : _T_1323) :
                _T_1323;	// sequencer-master.scala:321:24
      wire _T_1359 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1325 ? io_op_bits_base_vp_scalar : _T_1260) :
                _T_1326) : _T_1326;	// sequencer-master.scala:321:24
      wire _T_1360 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1327 ? io_op_bits_base_vp_pred : _T_1261) : _T_1328)
                : _T_1328;	// sequencer-master.scala:321:24
      wire [3:0] _T_1361 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1329 ? io_op_bits_base_vp_id : _T_1262) : _T_1330) :
                _T_1330;	// sequencer-master.scala:321:24
      wire _T_1362 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1332 ? io_op_bits_base_vp_scalar : _T_1264) :
                _T_1333) : _T_1333;	// sequencer-master.scala:321:24
      wire _T_1363 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1334 ? io_op_bits_base_vp_pred : _T_1265) : _T_1335)
                : _T_1335;	// sequencer-master.scala:321:24
      wire [3:0] _T_1364 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (&tail | _T_1336 ? io_op_bits_base_vp_id : _T_1266) : _T_1337) :
                _T_1337;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1365 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (&tail | _T_1339 ? io_op_bits_base_vp_scalar : _T_1268) :
                _T_1340) : _T_1340;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1366 = io_op_bits_active_vamo & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (&tail | _T_1341 ? io_op_bits_base_vp_pred : _T_1269) : _T_1342)
                : _T_1342;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1367 = io_op_bits_active_vamo ? ~_T_314 & (io_op_bits_base_vp_valid & _T_291 ?
                io_op_bits_base_vp_valid : ~_T_291 & ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ?
                io_op_bits_base_vp_valid : ~_T_4 & _T_1289)) : _T_1289;	// sequencer-master.scala:272:28, :321:24
      wire _T_1368 = io_op_bits_active_vamo ? ~_T_315 & (io_op_bits_base_vp_valid & _T_292 ?
                io_op_bits_base_vp_valid : ~_T_292 & ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ?
                io_op_bits_base_vp_valid : ~_T_5 & _T_1296)) : _T_1296;	// sequencer-master.scala:272:28, :321:24
      wire _T_1369 = io_op_bits_active_vamo ? ~_T_316 & (io_op_bits_base_vp_valid & _T_293 ?
                io_op_bits_base_vp_valid : ~_T_293 & ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ?
                io_op_bits_base_vp_valid : ~_T_6 & _T_1303)) : _T_1303;	// sequencer-master.scala:272:28, :321:24
      wire _T_1370 = io_op_bits_active_vamo ? ~_T_317 & (io_op_bits_base_vp_valid & _T_294 ?
                io_op_bits_base_vp_valid : ~_T_294 & ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ?
                io_op_bits_base_vp_valid : ~_T_7 & _T_1310)) : _T_1310;	// sequencer-master.scala:272:28, :321:24
      wire _T_1371 = io_op_bits_active_vamo ? ~_T_318 & (io_op_bits_base_vp_valid & _T_295 ?
                io_op_bits_base_vp_valid : ~_T_295 & ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ?
                io_op_bits_base_vp_valid : ~_T_8 & _T_1317)) : _T_1317;	// sequencer-master.scala:272:28, :321:24
      wire _T_1372 = io_op_bits_active_vamo ? ~_T_319 & (io_op_bits_base_vp_valid & _T_296 ?
                io_op_bits_base_vp_valid : ~_T_296 & ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ?
                io_op_bits_base_vp_valid : ~_T_9 & _T_1324)) : _T_1324;	// sequencer-master.scala:272:28, :321:24
      wire _T_1373 = io_op_bits_active_vamo ? ~_T_320 & (io_op_bits_base_vp_valid & _T_297 ?
                io_op_bits_base_vp_valid : ~_T_297 & ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ?
                io_op_bits_base_vp_valid : ~_T_10 & _T_1331)) : _T_1331;	// sequencer-master.scala:272:28, :321:24
      wire _T_1374 = io_op_bits_active_vamo ? ~(&_T_2) & (io_op_bits_base_vp_valid & &_T_1 ?
                io_op_bits_base_vp_valid : ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ?
                io_op_bits_base_vp_valid : ~(&tail) & _T_1338)) : _T_1338;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1375 = io_op_bits_active_vamo & (_T_314 | _T_291 | _T_132 | _T_4);	// sequencer-master.scala:289:23
      wire _T_1376 = io_op_bits_active_vamo & (_T_315 | _T_292 | _T_133 | _T_5);	// sequencer-master.scala:289:23
      wire _T_1377 = io_op_bits_active_vamo & (_T_316 | _T_293 | _T_134 | _T_6);	// sequencer-master.scala:289:23
      wire _T_1378 = io_op_bits_active_vamo & (_T_317 | _T_294 | _T_135 | _T_7);	// sequencer-master.scala:289:23
      wire _T_1379 = io_op_bits_active_vamo & (_T_318 | _T_295 | _T_136 | _T_8);	// sequencer-master.scala:289:23
      wire _T_1380 = io_op_bits_active_vamo & (_T_319 | _T_296 | _T_137 | _T_9);	// sequencer-master.scala:289:23
      wire _T_1381 = io_op_bits_active_vamo & (_T_320 | _T_297 | _T_138 | _T_10);	// sequencer-master.scala:289:23
      wire _T_1382 = io_op_bits_active_vamo & (&_T_2 | &_T_1 | &_T_0 | &tail);	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire _T_1383 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_314;	// sequencer-master.scala:363:24
      wire _T_1384 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_314 ? io_op_bits_base_vd_valid :
                ~_T_314 & ~_T_291 & ~_T_132 & ~_T_4 & _T_1270) : _T_1270;	// sequencer-master.scala:276:28, :363:24
      wire _T_1385 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_314;	// sequencer-master.scala:363:24
      wire _T_1386 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_314;	// sequencer-master.scala:363:24
      wire _T_1387 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_314;	// sequencer-master.scala:363:24
      wire _T_1388 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_315;	// sequencer-master.scala:363:24
      wire _T_1389 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_315 ? io_op_bits_base_vd_valid :
                ~_T_315 & ~_T_292 & ~_T_133 & ~_T_5 & _T_1271) : _T_1271;	// sequencer-master.scala:276:28, :363:24
      wire _T_1390 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_315;	// sequencer-master.scala:363:24
      wire _T_1391 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_315;	// sequencer-master.scala:363:24
      wire _T_1392 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_315;	// sequencer-master.scala:363:24
      wire _T_1393 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_316;	// sequencer-master.scala:363:24
      wire _T_1394 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_316 ? io_op_bits_base_vd_valid :
                ~_T_316 & ~_T_293 & ~_T_134 & ~_T_6 & _T_1272) : _T_1272;	// sequencer-master.scala:276:28, :363:24
      wire _T_1395 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_316;	// sequencer-master.scala:363:24
      wire _T_1396 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_316;	// sequencer-master.scala:363:24
      wire _T_1397 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_316;	// sequencer-master.scala:363:24
      wire _T_1398 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_317;	// sequencer-master.scala:363:24
      wire _T_1399 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_317 ? io_op_bits_base_vd_valid :
                ~_T_317 & ~_T_294 & ~_T_135 & ~_T_7 & _T_1273) : _T_1273;	// sequencer-master.scala:276:28, :363:24
      wire _T_1400 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_317;	// sequencer-master.scala:363:24
      wire _T_1401 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_317;	// sequencer-master.scala:363:24
      wire _T_1402 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_317;	// sequencer-master.scala:363:24
      wire _T_1403 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_318;	// sequencer-master.scala:363:24
      wire _T_1404 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_318 ? io_op_bits_base_vd_valid :
                ~_T_318 & ~_T_295 & ~_T_136 & ~_T_8 & _T_1274) : _T_1274;	// sequencer-master.scala:276:28, :363:24
      wire _T_1405 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_318;	// sequencer-master.scala:363:24
      wire _T_1406 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_318;	// sequencer-master.scala:363:24
      wire _T_1407 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_318;	// sequencer-master.scala:363:24
      wire _T_1408 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_319;	// sequencer-master.scala:363:24
      wire _T_1409 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_319 ? io_op_bits_base_vd_valid :
                ~_T_319 & ~_T_296 & ~_T_137 & ~_T_9 & _T_1275) : _T_1275;	// sequencer-master.scala:276:28, :363:24
      wire _T_1410 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_319;	// sequencer-master.scala:363:24
      wire _T_1411 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_319;	// sequencer-master.scala:363:24
      wire _T_1412 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_319;	// sequencer-master.scala:363:24
      wire _T_1413 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_320;	// sequencer-master.scala:363:24
      wire _T_1414 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & _T_320 ? io_op_bits_base_vd_valid :
                ~_T_320 & ~_T_297 & ~_T_138 & ~_T_10 & _T_1276) : _T_1276;	// sequencer-master.scala:276:28, :363:24
      wire _T_1415 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_320;	// sequencer-master.scala:363:24
      wire _T_1416 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_320;	// sequencer-master.scala:363:24
      wire _T_1417 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & _T_320;	// sequencer-master.scala:363:24
      wire _T_1418 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & &_T_2;	// sequencer-master.scala:267:35, :363:24
      wire _T_1419 = io_op_bits_active_vamo ? (io_op_bits_base_vd_valid & &_T_2 ? io_op_bits_base_vd_valid :
                ~(&_T_2) & ~(&_T_1) & ~(&_T_0) & ~(&tail) & _T_1277) : _T_1277;	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_1420 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & &_T_2;	// sequencer-master.scala:267:35, :363:24
      wire _T_1421 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & &_T_2;	// sequencer-master.scala:267:35, :363:24
      wire _T_1422 = io_op_bits_active_vamo & io_op_bits_base_vd_valid & &_T_2;	// sequencer-master.scala:267:35, :363:24
      wire _T_1423 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire [3:0] _T_1424 = _T_1423 ? io_op_bits_base_vp_id : _T_1343;	// sequencer-master.scala:321:24
      wire _T_1425 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1426 = _T_1425 ? io_op_bits_base_vp_scalar : _T_1344;	// sequencer-master.scala:321:24
      wire _T_1427 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1428 = _T_1427 ? io_op_bits_base_vp_pred : _T_1345;	// sequencer-master.scala:321:24
      wire _T_1429 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire [3:0] _T_1430 = _T_1429 ? io_op_bits_base_vp_id : _T_1346;	// sequencer-master.scala:321:24
      wire _T_1431 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1432 = _T_1431 ? io_op_bits_base_vp_scalar : _T_1347;	// sequencer-master.scala:321:24
      wire _T_1433 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1434 = _T_1433 ? io_op_bits_base_vp_pred : _T_1348;	// sequencer-master.scala:321:24
      wire _T_1435 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire [3:0] _T_1436 = _T_1435 ? io_op_bits_base_vp_id : _T_1349;	// sequencer-master.scala:321:24
      wire _T_1437 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1438 = _T_1437 ? io_op_bits_base_vp_scalar : _T_1350;	// sequencer-master.scala:321:24
      wire _T_1439 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1440 = _T_1439 ? io_op_bits_base_vp_pred : _T_1351;	// sequencer-master.scala:321:24
      wire _T_1441 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire [3:0] _T_1442 = _T_1441 ? io_op_bits_base_vp_id : _T_1352;	// sequencer-master.scala:321:24
      wire _T_1443 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1444 = _T_1443 ? io_op_bits_base_vp_scalar : _T_1353;	// sequencer-master.scala:321:24
      wire _T_1445 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1446 = _T_1445 ? io_op_bits_base_vp_pred : _T_1354;	// sequencer-master.scala:321:24
      wire _T_1447 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire [3:0] _T_1448 = _T_1447 ? io_op_bits_base_vp_id : _T_1355;	// sequencer-master.scala:321:24
      wire _T_1449 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1450 = _T_1449 ? io_op_bits_base_vp_scalar : _T_1356;	// sequencer-master.scala:321:24
      wire _T_1451 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1452 = _T_1451 ? io_op_bits_base_vp_pred : _T_1357;	// sequencer-master.scala:321:24
      wire _T_1453 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire [3:0] _T_1454 = _T_1453 ? io_op_bits_base_vp_id : _T_1358;	// sequencer-master.scala:321:24
      wire _T_1455 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1456 = _T_1455 ? io_op_bits_base_vp_scalar : _T_1359;	// sequencer-master.scala:321:24
      wire _T_1457 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1458 = _T_1457 ? io_op_bits_base_vp_pred : _T_1360;	// sequencer-master.scala:321:24
      wire _T_1459 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire [3:0] _T_1460 = _T_1459 ? io_op_bits_base_vp_id : _T_1361;	// sequencer-master.scala:321:24
      wire _T_1461 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1462 = _T_1461 ? io_op_bits_base_vp_scalar : _T_1362;	// sequencer-master.scala:321:24
      wire _T_1463 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1464 = _T_1463 ? io_op_bits_base_vp_pred : _T_1363;	// sequencer-master.scala:321:24
      wire _T_1465 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire [3:0] _T_1466 = _T_1465 ? io_op_bits_base_vp_id : _T_1364;	// sequencer-master.scala:321:24
      wire _T_1467 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1468 = _T_1467 ? io_op_bits_base_vp_scalar : _T_1365;	// sequencer-master.scala:321:24
      wire _T_1469 = io_op_bits_active_vldx & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1470 = _T_1469 ? io_op_bits_base_vp_pred : _T_1366;	// sequencer-master.scala:321:24
      wire _T_1471 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ?
                io_op_bits_base_vp_valid : ~_T_4 & _T_1367) : _T_1367;	// sequencer-master.scala:272:28, :321:24
      wire _T_1472 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ?
                io_op_bits_base_vp_valid : ~_T_5 & _T_1368) : _T_1368;	// sequencer-master.scala:272:28, :321:24
      wire _T_1473 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ?
                io_op_bits_base_vp_valid : ~_T_6 & _T_1369) : _T_1369;	// sequencer-master.scala:272:28, :321:24
      wire _T_1474 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ?
                io_op_bits_base_vp_valid : ~_T_7 & _T_1370) : _T_1370;	// sequencer-master.scala:272:28, :321:24
      wire _T_1475 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ?
                io_op_bits_base_vp_valid : ~_T_8 & _T_1371) : _T_1371;	// sequencer-master.scala:272:28, :321:24
      wire _T_1476 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ?
                io_op_bits_base_vp_valid : ~_T_9 & _T_1372) : _T_1372;	// sequencer-master.scala:272:28, :321:24
      wire _T_1477 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ?
                io_op_bits_base_vp_valid : ~_T_10 & _T_1373) : _T_1373;	// sequencer-master.scala:272:28, :321:24
      wire _T_1478 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ?
                io_op_bits_base_vp_valid : ~(&tail) & _T_1374) : _T_1374;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire [9:0] _T_1479 = io_op_bits_active_vldx ? (_T_291 | _T_132 | _T_4 | _T_1375 ? io_op_bits_fn_union : _T_1279)
                : _T_1375 ? io_op_bits_fn_union : _T_1279;	// sequencer-master.scala:289:23
      wire [9:0] _T_1480 = io_op_bits_active_vldx ? (_T_292 | _T_133 | _T_5 | _T_1376 ? io_op_bits_fn_union : _T_1280)
                : _T_1376 ? io_op_bits_fn_union : _T_1280;	// sequencer-master.scala:289:23
      wire [9:0] _T_1481 = io_op_bits_active_vldx ? (_T_293 | _T_134 | _T_6 | _T_1377 ? io_op_bits_fn_union : _T_1281)
                : _T_1377 ? io_op_bits_fn_union : _T_1281;	// sequencer-master.scala:289:23
      wire [9:0] _T_1482 = io_op_bits_active_vldx ? (_T_294 | _T_135 | _T_7 | _T_1378 ? io_op_bits_fn_union : _T_1282)
                : _T_1378 ? io_op_bits_fn_union : _T_1282;	// sequencer-master.scala:289:23
      wire [9:0] _T_1483 = io_op_bits_active_vldx ? (_T_295 | _T_136 | _T_8 | _T_1379 ? io_op_bits_fn_union : _T_1283)
                : _T_1379 ? io_op_bits_fn_union : _T_1283;	// sequencer-master.scala:289:23
      wire [9:0] _T_1484 = io_op_bits_active_vldx ? (_T_296 | _T_137 | _T_9 | _T_1380 ? io_op_bits_fn_union : _T_1284)
                : _T_1380 ? io_op_bits_fn_union : _T_1284;	// sequencer-master.scala:289:23
      wire [9:0] _T_1485 = io_op_bits_active_vldx ? (_T_297 | _T_138 | _T_10 | _T_1381 ? io_op_bits_fn_union :
                _T_1285) : _T_1381 ? io_op_bits_fn_union : _T_1285;	// sequencer-master.scala:289:23
      wire [9:0] _T_1486 = io_op_bits_active_vldx ? (&_T_1 | &_T_0 | &tail | _T_1382 ? io_op_bits_fn_union : _T_1286)
                : _T_1382 ? io_op_bits_fn_union : _T_1286;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire _T_1487 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_valid : ~_T_291 & ~_T_132 & ~_T_4 &
                _T_1384) : _T_1384);	// sequencer-master.scala:276:28, :363:24
      wire _T_1488 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_valid : ~_T_292 & ~_T_133 & ~_T_5 &
                _T_1389) : _T_1389);	// sequencer-master.scala:276:28, :363:24
      wire _T_1489 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_valid : ~_T_293 & ~_T_134 & ~_T_6 &
                _T_1394) : _T_1394);	// sequencer-master.scala:276:28, :363:24
      wire _T_1490 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_valid : ~_T_294 & ~_T_135 & ~_T_7 &
                _T_1399) : _T_1399);	// sequencer-master.scala:276:28, :363:24
      wire _T_1491 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_valid : ~_T_295 & ~_T_136 & ~_T_8 &
                _T_1404) : _T_1404);	// sequencer-master.scala:276:28, :363:24
      wire _T_1492 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_valid : ~_T_296 & ~_T_137 & ~_T_9 &
                _T_1409) : _T_1409);	// sequencer-master.scala:276:28, :363:24
      wire _T_1493 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_valid : ~_T_297 & ~_T_138 & ~_T_10
                & _T_1414) : _T_1414);	// sequencer-master.scala:276:28, :363:24
      wire _T_1494 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_valid : ~(&_T_1) & ~(&_T_0) &
                ~(&tail) & _T_1419) : _T_1419);	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      wire _T_1495 = io_op_bits_active_vstx & (_T_291 | _T_132 | _T_4);	// sequencer-master.scala:289:23
      wire _T_1496 = io_op_bits_active_vstx & (_T_292 | _T_133 | _T_5);	// sequencer-master.scala:289:23
      wire _T_1497 = io_op_bits_active_vstx & (_T_293 | _T_134 | _T_6);	// sequencer-master.scala:289:23
      wire _T_1498 = io_op_bits_active_vstx & (_T_294 | _T_135 | _T_7);	// sequencer-master.scala:289:23
      wire _T_1499 = io_op_bits_active_vstx & (_T_295 | _T_136 | _T_8);	// sequencer-master.scala:289:23
      wire _T_1500 = io_op_bits_active_vstx & (_T_296 | _T_137 | _T_9);	// sequencer-master.scala:289:23
      wire _T_1501 = io_op_bits_active_vstx & (_T_297 | _T_138 | _T_10);	// sequencer-master.scala:289:23
      wire _T_1502 = io_op_bits_active_vstx & (&_T_1 | &_T_0 | &tail);	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      wire [3:0] _T_1503 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1423 ? io_op_bits_base_vp_id : _T_1343) : _T_1424) :
                _T_1424;	// sequencer-master.scala:321:24
      wire _T_1504 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_291 ? io_op_bits_base_vp_valid :
                ~_T_291 & ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid : ~_T_4 &
                _T_1471)) : _T_1471;	// sequencer-master.scala:272:28, :321:24
      wire _T_1505 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1425 ? io_op_bits_base_vp_scalar : _T_1344) :
                _T_1426) : _T_1426;	// sequencer-master.scala:321:24
      wire _T_1506 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_4 | _T_1427 ? io_op_bits_base_vp_pred : _T_1345) : _T_1428)
                : _T_1428;	// sequencer-master.scala:321:24
      wire [3:0] _T_1507 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1429 ? io_op_bits_base_vp_id : _T_1346) : _T_1430) :
                _T_1430;	// sequencer-master.scala:321:24
      wire _T_1508 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_292 ? io_op_bits_base_vp_valid :
                ~_T_292 & ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid : ~_T_5 &
                _T_1472)) : _T_1472;	// sequencer-master.scala:272:28, :321:24
      wire _T_1509 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1431 ? io_op_bits_base_vp_scalar : _T_1347) :
                _T_1432) : _T_1432;	// sequencer-master.scala:321:24
      wire _T_1510 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_5 | _T_1433 ? io_op_bits_base_vp_pred : _T_1348) : _T_1434)
                : _T_1434;	// sequencer-master.scala:321:24
      wire [3:0] _T_1511 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1435 ? io_op_bits_base_vp_id : _T_1349) : _T_1436) :
                _T_1436;	// sequencer-master.scala:321:24
      wire _T_1512 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_293 ? io_op_bits_base_vp_valid :
                ~_T_293 & ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid : ~_T_6 &
                _T_1473)) : _T_1473;	// sequencer-master.scala:272:28, :321:24
      wire _T_1513 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1437 ? io_op_bits_base_vp_scalar : _T_1350) :
                _T_1438) : _T_1438;	// sequencer-master.scala:321:24
      wire _T_1514 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_6 | _T_1439 ? io_op_bits_base_vp_pred : _T_1351) : _T_1440)
                : _T_1440;	// sequencer-master.scala:321:24
      wire [3:0] _T_1515 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1441 ? io_op_bits_base_vp_id : _T_1352) : _T_1442) :
                _T_1442;	// sequencer-master.scala:321:24
      wire _T_1516 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_294 ? io_op_bits_base_vp_valid :
                ~_T_294 & ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid : ~_T_7 &
                _T_1474)) : _T_1474;	// sequencer-master.scala:272:28, :321:24
      wire _T_1517 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1443 ? io_op_bits_base_vp_scalar : _T_1353) :
                _T_1444) : _T_1444;	// sequencer-master.scala:321:24
      wire _T_1518 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_7 | _T_1445 ? io_op_bits_base_vp_pred : _T_1354) : _T_1446)
                : _T_1446;	// sequencer-master.scala:321:24
      wire [3:0] _T_1519 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1447 ? io_op_bits_base_vp_id : _T_1355) : _T_1448) :
                _T_1448;	// sequencer-master.scala:321:24
      wire _T_1520 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_295 ? io_op_bits_base_vp_valid :
                ~_T_295 & ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid : ~_T_8 &
                _T_1475)) : _T_1475;	// sequencer-master.scala:272:28, :321:24
      wire _T_1521 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1449 ? io_op_bits_base_vp_scalar : _T_1356) :
                _T_1450) : _T_1450;	// sequencer-master.scala:321:24
      wire _T_1522 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_8 | _T_1451 ? io_op_bits_base_vp_pred : _T_1357) : _T_1452)
                : _T_1452;	// sequencer-master.scala:321:24
      wire [3:0] _T_1523 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1453 ? io_op_bits_base_vp_id : _T_1358) : _T_1454) :
                _T_1454;	// sequencer-master.scala:321:24
      wire _T_1524 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_296 ? io_op_bits_base_vp_valid :
                ~_T_296 & ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid : ~_T_9 &
                _T_1476)) : _T_1476;	// sequencer-master.scala:272:28, :321:24
      wire _T_1525 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1455 ? io_op_bits_base_vp_scalar : _T_1359) :
                _T_1456) : _T_1456;	// sequencer-master.scala:321:24
      wire _T_1526 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_9 | _T_1457 ? io_op_bits_base_vp_pred : _T_1360) : _T_1458)
                : _T_1458;	// sequencer-master.scala:321:24
      wire [3:0] _T_1527 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1459 ? io_op_bits_base_vp_id : _T_1361) : _T_1460) :
                _T_1460;	// sequencer-master.scala:321:24
      wire _T_1528 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & _T_297 ? io_op_bits_base_vp_valid :
                ~_T_297 & ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid : ~_T_10 &
                _T_1477)) : _T_1477;	// sequencer-master.scala:272:28, :321:24
      wire _T_1529 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1461 ? io_op_bits_base_vp_scalar : _T_1362) :
                _T_1462) : _T_1462;	// sequencer-master.scala:321:24
      wire _T_1530 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (_T_10 | _T_1463 ? io_op_bits_base_vp_pred : _T_1363) : _T_1464)
                : _T_1464;	// sequencer-master.scala:321:24
      wire [3:0] _T_1531 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_id :
                io_op_bits_base_vp_valid ? (&tail | _T_1465 ? io_op_bits_base_vp_id : _T_1364) : _T_1466) :
                _T_1466;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1532 = io_op_bits_active_vstx ? (io_op_bits_base_vp_valid & &_T_1 ? io_op_bits_base_vp_valid :
                ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                ~(&tail) & _T_1478)) : _T_1478;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1533 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_scalar :
                io_op_bits_base_vp_valid ? (&tail | _T_1467 ? io_op_bits_base_vp_scalar : _T_1365) :
                _T_1468) : _T_1468;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1534 = io_op_bits_active_vstx & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_pred :
                io_op_bits_base_vp_valid ? (&tail | _T_1469 ? io_op_bits_base_vp_pred : _T_1366) : _T_1470)
                : _T_1470;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1535 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire [3:0] _T_1536 = _T_1535 ? io_op_bits_base_vp_id : _T_1503;	// sequencer-master.scala:321:24
      wire _T_1537 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1538 = _T_1537 ? io_op_bits_base_vp_scalar : _T_1505;	// sequencer-master.scala:321:24
      wire _T_1539 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_4;	// sequencer-master.scala:321:24
      wire _T_1540 = _T_1539 ? io_op_bits_base_vp_pred : _T_1506;	// sequencer-master.scala:321:24
      wire _T_1541 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire [3:0] _T_1542 = _T_1541 ? io_op_bits_base_vp_id : _T_1507;	// sequencer-master.scala:321:24
      wire _T_1543 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1544 = _T_1543 ? io_op_bits_base_vp_scalar : _T_1509;	// sequencer-master.scala:321:24
      wire _T_1545 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_5;	// sequencer-master.scala:321:24
      wire _T_1546 = _T_1545 ? io_op_bits_base_vp_pred : _T_1510;	// sequencer-master.scala:321:24
      wire _T_1547 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire [3:0] _T_1548 = _T_1547 ? io_op_bits_base_vp_id : _T_1511;	// sequencer-master.scala:321:24
      wire _T_1549 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1550 = _T_1549 ? io_op_bits_base_vp_scalar : _T_1513;	// sequencer-master.scala:321:24
      wire _T_1551 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_6;	// sequencer-master.scala:321:24
      wire _T_1552 = _T_1551 ? io_op_bits_base_vp_pred : _T_1514;	// sequencer-master.scala:321:24
      wire _T_1553 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire [3:0] _T_1554 = _T_1553 ? io_op_bits_base_vp_id : _T_1515;	// sequencer-master.scala:321:24
      wire _T_1555 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1556 = _T_1555 ? io_op_bits_base_vp_scalar : _T_1517;	// sequencer-master.scala:321:24
      wire _T_1557 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_7;	// sequencer-master.scala:321:24
      wire _T_1558 = _T_1557 ? io_op_bits_base_vp_pred : _T_1518;	// sequencer-master.scala:321:24
      wire _T_1559 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire [3:0] _T_1560 = _T_1559 ? io_op_bits_base_vp_id : _T_1519;	// sequencer-master.scala:321:24
      wire _T_1561 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1562 = _T_1561 ? io_op_bits_base_vp_scalar : _T_1521;	// sequencer-master.scala:321:24
      wire _T_1563 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_8;	// sequencer-master.scala:321:24
      wire _T_1564 = _T_1563 ? io_op_bits_base_vp_pred : _T_1522;	// sequencer-master.scala:321:24
      wire _T_1565 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire [3:0] _T_1566 = _T_1565 ? io_op_bits_base_vp_id : _T_1523;	// sequencer-master.scala:321:24
      wire _T_1567 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1568 = _T_1567 ? io_op_bits_base_vp_scalar : _T_1525;	// sequencer-master.scala:321:24
      wire _T_1569 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_9;	// sequencer-master.scala:321:24
      wire _T_1570 = _T_1569 ? io_op_bits_base_vp_pred : _T_1526;	// sequencer-master.scala:321:24
      wire _T_1571 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire [3:0] _T_1572 = _T_1571 ? io_op_bits_base_vp_id : _T_1527;	// sequencer-master.scala:321:24
      wire _T_1573 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1574 = _T_1573 ? io_op_bits_base_vp_scalar : _T_1529;	// sequencer-master.scala:321:24
      wire _T_1575 = io_op_bits_active_vld & io_op_bits_base_vp_valid & _T_10;	// sequencer-master.scala:321:24
      wire _T_1576 = _T_1575 ? io_op_bits_base_vp_pred : _T_1530;	// sequencer-master.scala:321:24
      wire _T_1577 = io_op_bits_active_vld & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire [3:0] _T_1578 = _T_1577 ? io_op_bits_base_vp_id : _T_1531;	// sequencer-master.scala:321:24
      wire _T_1579 = io_op_bits_active_vld & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1580 = _T_1579 ? io_op_bits_base_vp_scalar : _T_1533;	// sequencer-master.scala:321:24
      wire _T_1581 = io_op_bits_active_vld & io_op_bits_base_vp_valid & &tail;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      wire _T_1582 = _T_1581 ? io_op_bits_base_vp_pred : _T_1534;	// sequencer-master.scala:321:24
      wire _T_1583 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ?
                io_op_bits_base_vp_valid : ~_T_4 & _T_1504) : _T_1504;	// sequencer-master.scala:272:28, :321:24
      wire _T_1584 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ?
                io_op_bits_base_vp_valid : ~_T_5 & _T_1508) : _T_1508;	// sequencer-master.scala:272:28, :321:24
      wire _T_1585 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ?
                io_op_bits_base_vp_valid : ~_T_6 & _T_1512) : _T_1512;	// sequencer-master.scala:272:28, :321:24
      wire _T_1586 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ?
                io_op_bits_base_vp_valid : ~_T_7 & _T_1516) : _T_1516;	// sequencer-master.scala:272:28, :321:24
      wire _T_1587 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ?
                io_op_bits_base_vp_valid : ~_T_8 & _T_1520) : _T_1520;	// sequencer-master.scala:272:28, :321:24
      wire _T_1588 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ?
                io_op_bits_base_vp_valid : ~_T_9 & _T_1524) : _T_1524;	// sequencer-master.scala:272:28, :321:24
      wire _T_1589 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ?
                io_op_bits_base_vp_valid : ~_T_10 & _T_1528) : _T_1528;	// sequencer-master.scala:272:28, :321:24
      wire _T_1590 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ?
                io_op_bits_base_vp_valid : ~(&tail) & _T_1532) : _T_1532;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      wire _T_1591 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1592 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & e_0_base_vs1_valid) : e_0_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1593 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1594 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1595 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1596 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1597 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & e_1_base_vs1_valid) : e_1_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1598 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1599 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1600 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1601 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1602 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & e_2_base_vs1_valid) : e_2_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1603 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1604 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1605 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1606 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1607 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & e_3_base_vs1_valid) : e_3_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1608 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1609 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1610 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1611 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1612 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & e_4_base_vs1_valid) : e_4_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1613 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1614 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1615 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1616 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1617 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & e_5_base_vs1_valid) : e_5_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1618 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1619 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1620 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1621 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1622 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid :
                ~_T_10 & e_6_base_vs1_valid) : e_6_base_vs1_valid;	// sequencer-master.scala:136:44, :273:29, :329:29
      wire _T_1623 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1624 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1625 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1626 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1627 = io_op_bits_active_vint ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid :
                ~(&tail) & e_7_base_vs1_valid) : e_7_base_vs1_valid;	// sequencer-master.scala:136:44, :267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1628 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1629 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1630 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1631 = io_op_bits_active_vint & _T_4;	// sequencer-master.scala:230:21
      wire _T_1632 = io_op_bits_active_vint & _T_5;	// sequencer-master.scala:230:21
      wire _T_1633 = io_op_bits_active_vint & _T_6;	// sequencer-master.scala:230:21
      wire _T_1634 = io_op_bits_active_vint & _T_7;	// sequencer-master.scala:230:21
      wire _T_1635 = io_op_bits_active_vint & _T_8;	// sequencer-master.scala:230:21
      wire _T_1636 = io_op_bits_active_vint & _T_9;	// sequencer-master.scala:230:21
      wire _T_1637 = io_op_bits_active_vint & _T_10;	// sequencer-master.scala:230:21
      wire _T_1638 = io_op_bits_active_vint & &tail;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [7:0] _T_1639 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_4 | _T_1591 ?
                io_op_bits_base_vs1_id : e_0_base_vs1_id) : _T_1591 ? io_op_bits_base_vs1_id :
                e_0_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1640 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & _T_1592) : _T_1592;	// sequencer-master.scala:273:29, :329:29
      wire _T_1641 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_4 | _T_1593 ?
                io_op_bits_base_vs1_scalar : e_0_base_vs1_scalar) : _T_1593 ? io_op_bits_base_vs1_scalar :
                e_0_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1642 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_4 | _T_1594 ?
                io_op_bits_base_vs1_pred : e_0_base_vs1_pred) : _T_1594 ? io_op_bits_base_vs1_pred :
                e_0_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1643 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_4 | _T_1595 ?
                io_op_bits_base_vs1_prec : e_0_base_vs1_prec) : _T_1595 ? io_op_bits_base_vs1_prec :
                e_0_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1644 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_5 | _T_1596 ?
                io_op_bits_base_vs1_id : e_1_base_vs1_id) : _T_1596 ? io_op_bits_base_vs1_id :
                e_1_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1645 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & _T_1597) : _T_1597;	// sequencer-master.scala:273:29, :329:29
      wire _T_1646 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_5 | _T_1598 ?
                io_op_bits_base_vs1_scalar : e_1_base_vs1_scalar) : _T_1598 ? io_op_bits_base_vs1_scalar :
                e_1_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1647 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_5 | _T_1599 ?
                io_op_bits_base_vs1_pred : e_1_base_vs1_pred) : _T_1599 ? io_op_bits_base_vs1_pred :
                e_1_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1648 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_5 | _T_1600 ?
                io_op_bits_base_vs1_prec : e_1_base_vs1_prec) : _T_1600 ? io_op_bits_base_vs1_prec :
                e_1_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1649 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_6 | _T_1601 ?
                io_op_bits_base_vs1_id : e_2_base_vs1_id) : _T_1601 ? io_op_bits_base_vs1_id :
                e_2_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1650 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & _T_1602) : _T_1602;	// sequencer-master.scala:273:29, :329:29
      wire _T_1651 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_6 | _T_1603 ?
                io_op_bits_base_vs1_scalar : e_2_base_vs1_scalar) : _T_1603 ? io_op_bits_base_vs1_scalar :
                e_2_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1652 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_6 | _T_1604 ?
                io_op_bits_base_vs1_pred : e_2_base_vs1_pred) : _T_1604 ? io_op_bits_base_vs1_pred :
                e_2_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1653 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_6 | _T_1605 ?
                io_op_bits_base_vs1_prec : e_2_base_vs1_prec) : _T_1605 ? io_op_bits_base_vs1_prec :
                e_2_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1654 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_7 | _T_1606 ?
                io_op_bits_base_vs1_id : e_3_base_vs1_id) : _T_1606 ? io_op_bits_base_vs1_id :
                e_3_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1655 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & _T_1607) : _T_1607;	// sequencer-master.scala:273:29, :329:29
      wire _T_1656 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_7 | _T_1608 ?
                io_op_bits_base_vs1_scalar : e_3_base_vs1_scalar) : _T_1608 ? io_op_bits_base_vs1_scalar :
                e_3_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1657 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_7 | _T_1609 ?
                io_op_bits_base_vs1_pred : e_3_base_vs1_pred) : _T_1609 ? io_op_bits_base_vs1_pred :
                e_3_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1658 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_7 | _T_1610 ?
                io_op_bits_base_vs1_prec : e_3_base_vs1_prec) : _T_1610 ? io_op_bits_base_vs1_prec :
                e_3_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1659 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_8 | _T_1611 ?
                io_op_bits_base_vs1_id : e_4_base_vs1_id) : _T_1611 ? io_op_bits_base_vs1_id :
                e_4_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1660 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & _T_1612) : _T_1612;	// sequencer-master.scala:273:29, :329:29
      wire _T_1661 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_8 | _T_1613 ?
                io_op_bits_base_vs1_scalar : e_4_base_vs1_scalar) : _T_1613 ? io_op_bits_base_vs1_scalar :
                e_4_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1662 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_8 | _T_1614 ?
                io_op_bits_base_vs1_pred : e_4_base_vs1_pred) : _T_1614 ? io_op_bits_base_vs1_pred :
                e_4_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1663 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_8 | _T_1615 ?
                io_op_bits_base_vs1_prec : e_4_base_vs1_prec) : _T_1615 ? io_op_bits_base_vs1_prec :
                e_4_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1664 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_9 | _T_1616 ?
                io_op_bits_base_vs1_id : e_5_base_vs1_id) : _T_1616 ? io_op_bits_base_vs1_id :
                e_5_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1665 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & _T_1617) : _T_1617;	// sequencer-master.scala:273:29, :329:29
      wire _T_1666 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_9 | _T_1618 ?
                io_op_bits_base_vs1_scalar : e_5_base_vs1_scalar) : _T_1618 ? io_op_bits_base_vs1_scalar :
                e_5_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1667 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_9 | _T_1619 ?
                io_op_bits_base_vs1_pred : e_5_base_vs1_pred) : _T_1619 ? io_op_bits_base_vs1_pred :
                e_5_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1668 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_9 | _T_1620 ?
                io_op_bits_base_vs1_prec : e_5_base_vs1_prec) : _T_1620 ? io_op_bits_base_vs1_prec :
                e_5_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1669 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_10 | _T_1621 ?
                io_op_bits_base_vs1_id : e_6_base_vs1_id) : _T_1621 ? io_op_bits_base_vs1_id :
                e_6_base_vs1_id;	// sequencer-master.scala:141:29, :329:29
      wire _T_1670 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid :
                ~_T_10 & _T_1622) : _T_1622;	// sequencer-master.scala:273:29, :329:29
      wire _T_1671 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_10 | _T_1623 ?
                io_op_bits_base_vs1_scalar : e_6_base_vs1_scalar) : _T_1623 ? io_op_bits_base_vs1_scalar :
                e_6_base_vs1_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      wire _T_1672 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_10 | _T_1624 ?
                io_op_bits_base_vs1_pred : e_6_base_vs1_pred) : _T_1624 ? io_op_bits_base_vs1_pred :
                e_6_base_vs1_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      wire [1:0] _T_1673 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (_T_10 | _T_1625 ?
                io_op_bits_base_vs1_prec : e_6_base_vs1_prec) : _T_1625 ? io_op_bits_base_vs1_prec :
                e_6_base_vs1_prec;	// sequencer-master.scala:329:29
      wire [7:0] _T_1674 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (&tail | _T_1626 ?
                io_op_bits_base_vs1_id : e_7_base_vs1_id) : _T_1626 ? io_op_bits_base_vs1_id :
                e_7_base_vs1_id;	// sequencer-master.scala:141:29, :267:35, :329:29, util.scala:94:11
      wire _T_1675 = io_op_bits_active_vipred ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid :
                ~(&tail) & _T_1627) : _T_1627;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1676 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (&tail | _T_1628 ?
                io_op_bits_base_vs1_scalar : e_7_base_vs1_scalar) : _T_1628 ? io_op_bits_base_vs1_scalar :
                e_7_base_vs1_scalar;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:37, util.scala:94:11
      wire _T_1677 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (&tail | _T_1629 ?
                io_op_bits_base_vs1_pred : e_7_base_vs1_pred) : _T_1629 ? io_op_bits_base_vs1_pred :
                e_7_base_vs1_pred;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:31, util.scala:94:11
      wire [1:0] _T_1678 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid ? (&tail | _T_1630 ?
                io_op_bits_base_vs1_prec : e_7_base_vs1_prec) : _T_1630 ? io_op_bits_base_vs1_prec :
                e_7_base_vs1_prec;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1679 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1680 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & _T_1640) : _T_1640;	// sequencer-master.scala:273:29, :329:29
      wire _T_1681 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1682 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1683 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1684 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1685 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & _T_1645) : _T_1645;	// sequencer-master.scala:273:29, :329:29
      wire _T_1686 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1687 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1688 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1689 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1690 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & _T_1650) : _T_1650;	// sequencer-master.scala:273:29, :329:29
      wire _T_1691 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1692 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1693 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1694 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1695 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & _T_1655) : _T_1655;	// sequencer-master.scala:273:29, :329:29
      wire _T_1696 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1697 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1698 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1699 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1700 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & _T_1660) : _T_1660;	// sequencer-master.scala:273:29, :329:29
      wire _T_1701 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1702 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1703 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1704 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1705 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & _T_1665) : _T_1665;	// sequencer-master.scala:273:29, :329:29
      wire _T_1706 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1707 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1708 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1709 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1710 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid :
                ~_T_10 & _T_1670) : _T_1670;	// sequencer-master.scala:273:29, :329:29
      wire _T_1711 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1712 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1713 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1714 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1715 = io_op_bits_active_vimul ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid :
                ~(&tail) & _T_1675) : _T_1675;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1716 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1717 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1718 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1719 = io_op_bits_active_vimul & _T_4;	// sequencer-master.scala:230:21
      wire _T_1720 = io_op_bits_active_vimul & _T_5;	// sequencer-master.scala:230:21
      wire _T_1721 = io_op_bits_active_vimul & _T_6;	// sequencer-master.scala:230:21
      wire _T_1722 = io_op_bits_active_vimul & _T_7;	// sequencer-master.scala:230:21
      wire _T_1723 = io_op_bits_active_vimul & _T_8;	// sequencer-master.scala:230:21
      wire _T_1724 = io_op_bits_active_vimul & _T_9;	// sequencer-master.scala:230:21
      wire _T_1725 = io_op_bits_active_vimul & _T_10;	// sequencer-master.scala:230:21
      wire _T_1726 = io_op_bits_active_vimul & &tail;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [7:0] _T_1727 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1679 ?
                io_op_bits_base_vs1_id : _T_1639) : _T_1679 ? io_op_bits_base_vs1_id : _T_1639;	// sequencer-master.scala:329:29
      wire _T_1728 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1681 ?
                io_op_bits_base_vs1_scalar : _T_1641) : _T_1681 ? io_op_bits_base_vs1_scalar : _T_1641;	// sequencer-master.scala:329:29
      wire _T_1729 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1682 ?
                io_op_bits_base_vs1_pred : _T_1642) : _T_1682 ? io_op_bits_base_vs1_pred : _T_1642;	// sequencer-master.scala:329:29
      wire [1:0] _T_1730 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1683 ?
                io_op_bits_base_vs1_prec : _T_1643) : _T_1683 ? io_op_bits_base_vs1_prec : _T_1643;	// sequencer-master.scala:329:29
      wire [7:0] _T_1731 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1684 ?
                io_op_bits_base_vs1_id : _T_1644) : _T_1684 ? io_op_bits_base_vs1_id : _T_1644;	// sequencer-master.scala:329:29
      wire _T_1732 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1686 ?
                io_op_bits_base_vs1_scalar : _T_1646) : _T_1686 ? io_op_bits_base_vs1_scalar : _T_1646;	// sequencer-master.scala:329:29
      wire _T_1733 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1687 ?
                io_op_bits_base_vs1_pred : _T_1647) : _T_1687 ? io_op_bits_base_vs1_pred : _T_1647;	// sequencer-master.scala:329:29
      wire [1:0] _T_1734 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1688 ?
                io_op_bits_base_vs1_prec : _T_1648) : _T_1688 ? io_op_bits_base_vs1_prec : _T_1648;	// sequencer-master.scala:329:29
      wire [7:0] _T_1735 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1689 ?
                io_op_bits_base_vs1_id : _T_1649) : _T_1689 ? io_op_bits_base_vs1_id : _T_1649;	// sequencer-master.scala:329:29
      wire _T_1736 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1691 ?
                io_op_bits_base_vs1_scalar : _T_1651) : _T_1691 ? io_op_bits_base_vs1_scalar : _T_1651;	// sequencer-master.scala:329:29
      wire _T_1737 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1692 ?
                io_op_bits_base_vs1_pred : _T_1652) : _T_1692 ? io_op_bits_base_vs1_pred : _T_1652;	// sequencer-master.scala:329:29
      wire [1:0] _T_1738 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1693 ?
                io_op_bits_base_vs1_prec : _T_1653) : _T_1693 ? io_op_bits_base_vs1_prec : _T_1653;	// sequencer-master.scala:329:29
      wire [7:0] _T_1739 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1694 ?
                io_op_bits_base_vs1_id : _T_1654) : _T_1694 ? io_op_bits_base_vs1_id : _T_1654;	// sequencer-master.scala:329:29
      wire _T_1740 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1696 ?
                io_op_bits_base_vs1_scalar : _T_1656) : _T_1696 ? io_op_bits_base_vs1_scalar : _T_1656;	// sequencer-master.scala:329:29
      wire _T_1741 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1697 ?
                io_op_bits_base_vs1_pred : _T_1657) : _T_1697 ? io_op_bits_base_vs1_pred : _T_1657;	// sequencer-master.scala:329:29
      wire [1:0] _T_1742 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1698 ?
                io_op_bits_base_vs1_prec : _T_1658) : _T_1698 ? io_op_bits_base_vs1_prec : _T_1658;	// sequencer-master.scala:329:29
      wire [7:0] _T_1743 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1699 ?
                io_op_bits_base_vs1_id : _T_1659) : _T_1699 ? io_op_bits_base_vs1_id : _T_1659;	// sequencer-master.scala:329:29
      wire _T_1744 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1701 ?
                io_op_bits_base_vs1_scalar : _T_1661) : _T_1701 ? io_op_bits_base_vs1_scalar : _T_1661;	// sequencer-master.scala:329:29
      wire _T_1745 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1702 ?
                io_op_bits_base_vs1_pred : _T_1662) : _T_1702 ? io_op_bits_base_vs1_pred : _T_1662;	// sequencer-master.scala:329:29
      wire [1:0] _T_1746 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1703 ?
                io_op_bits_base_vs1_prec : _T_1663) : _T_1703 ? io_op_bits_base_vs1_prec : _T_1663;	// sequencer-master.scala:329:29
      wire [7:0] _T_1747 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1704 ?
                io_op_bits_base_vs1_id : _T_1664) : _T_1704 ? io_op_bits_base_vs1_id : _T_1664;	// sequencer-master.scala:329:29
      wire _T_1748 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1706 ?
                io_op_bits_base_vs1_scalar : _T_1666) : _T_1706 ? io_op_bits_base_vs1_scalar : _T_1666;	// sequencer-master.scala:329:29
      wire _T_1749 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1707 ?
                io_op_bits_base_vs1_pred : _T_1667) : _T_1707 ? io_op_bits_base_vs1_pred : _T_1667;	// sequencer-master.scala:329:29
      wire [1:0] _T_1750 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1708 ?
                io_op_bits_base_vs1_prec : _T_1668) : _T_1708 ? io_op_bits_base_vs1_prec : _T_1668;	// sequencer-master.scala:329:29
      wire [7:0] _T_1751 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1709 ?
                io_op_bits_base_vs1_id : _T_1669) : _T_1709 ? io_op_bits_base_vs1_id : _T_1669;	// sequencer-master.scala:329:29
      wire _T_1752 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1711 ?
                io_op_bits_base_vs1_scalar : _T_1671) : _T_1711 ? io_op_bits_base_vs1_scalar : _T_1671;	// sequencer-master.scala:329:29
      wire _T_1753 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1712 ?
                io_op_bits_base_vs1_pred : _T_1672) : _T_1712 ? io_op_bits_base_vs1_pred : _T_1672;	// sequencer-master.scala:329:29
      wire [1:0] _T_1754 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1713 ?
                io_op_bits_base_vs1_prec : _T_1673) : _T_1713 ? io_op_bits_base_vs1_prec : _T_1673;	// sequencer-master.scala:329:29
      wire [7:0] _T_1755 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (&tail | _T_1714 ?
                io_op_bits_base_vs1_id : _T_1674) : _T_1714 ? io_op_bits_base_vs1_id : _T_1674;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1756 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (&tail | _T_1716 ?
                io_op_bits_base_vs1_scalar : _T_1676) : _T_1716 ? io_op_bits_base_vs1_scalar : _T_1676;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1757 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (&tail | _T_1717 ?
                io_op_bits_base_vs1_pred : _T_1677) : _T_1717 ? io_op_bits_base_vs1_pred : _T_1677;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_1758 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid ? (&tail | _T_1718 ?
                io_op_bits_base_vs1_prec : _T_1678) : _T_1718 ? io_op_bits_base_vs1_prec : _T_1678;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1759 = io_op_bits_active_vidiv ? ~_T_132 & (io_op_bits_base_vs1_valid & _T_4 ?
                io_op_bits_base_vs1_valid : ~_T_4 & _T_1680) : _T_1680;	// sequencer-master.scala:273:29, :329:29
      wire _T_1760 = io_op_bits_active_vidiv ? ~_T_133 & (io_op_bits_base_vs1_valid & _T_5 ?
                io_op_bits_base_vs1_valid : ~_T_5 & _T_1685) : _T_1685;	// sequencer-master.scala:273:29, :329:29
      wire _T_1761 = io_op_bits_active_vidiv ? ~_T_134 & (io_op_bits_base_vs1_valid & _T_6 ?
                io_op_bits_base_vs1_valid : ~_T_6 & _T_1690) : _T_1690;	// sequencer-master.scala:273:29, :329:29
      wire _T_1762 = io_op_bits_active_vidiv ? ~_T_135 & (io_op_bits_base_vs1_valid & _T_7 ?
                io_op_bits_base_vs1_valid : ~_T_7 & _T_1695) : _T_1695;	// sequencer-master.scala:273:29, :329:29
      wire _T_1763 = io_op_bits_active_vidiv ? ~_T_136 & (io_op_bits_base_vs1_valid & _T_8 ?
                io_op_bits_base_vs1_valid : ~_T_8 & _T_1700) : _T_1700;	// sequencer-master.scala:273:29, :329:29
      wire _T_1764 = io_op_bits_active_vidiv ? ~_T_137 & (io_op_bits_base_vs1_valid & _T_9 ?
                io_op_bits_base_vs1_valid : ~_T_9 & _T_1705) : _T_1705;	// sequencer-master.scala:273:29, :329:29
      wire _T_1765 = io_op_bits_active_vidiv ? ~_T_138 & (io_op_bits_base_vs1_valid & _T_10 ?
                io_op_bits_base_vs1_valid : ~_T_10 & _T_1710) : _T_1710;	// sequencer-master.scala:273:29, :329:29
      wire _T_1766 = io_op_bits_active_vidiv ? ~(&_T_0) & (io_op_bits_base_vs1_valid & &tail ?
                io_op_bits_base_vs1_valid : ~(&tail) & _T_1715) : _T_1715;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1767 = io_op_bits_active_vidiv & (_T_132 | _T_4);	// sequencer-master.scala:231:25
      wire _T_1768 = io_op_bits_active_vidiv & (_T_133 | _T_5);	// sequencer-master.scala:231:25
      wire _T_1769 = io_op_bits_active_vidiv & (_T_134 | _T_6);	// sequencer-master.scala:231:25
      wire _T_1770 = io_op_bits_active_vidiv & (_T_135 | _T_7);	// sequencer-master.scala:231:25
      wire _T_1771 = io_op_bits_active_vidiv & (_T_136 | _T_8);	// sequencer-master.scala:231:25
      wire _T_1772 = io_op_bits_active_vidiv & (_T_137 | _T_9);	// sequencer-master.scala:231:25
      wire _T_1773 = io_op_bits_active_vidiv & (_T_138 | _T_10);	// sequencer-master.scala:231:25
      wire _T_1774 = io_op_bits_active_vidiv & (&_T_0 | &tail);	// sequencer-master.scala:231:25, :267:35, util.scala:94:11
      wire _T_1775 = io_op_bits_active_vidiv & (_T_132 | _T_4);	// sequencer-master.scala:232:25
      wire _T_1776 = io_op_bits_active_vidiv & (_T_133 | _T_5);	// sequencer-master.scala:232:25
      wire _T_1777 = io_op_bits_active_vidiv & (_T_134 | _T_6);	// sequencer-master.scala:232:25
      wire _T_1778 = io_op_bits_active_vidiv & (_T_135 | _T_7);	// sequencer-master.scala:232:25
      wire _T_1779 = io_op_bits_active_vidiv & (_T_136 | _T_8);	// sequencer-master.scala:232:25
      wire _T_1780 = io_op_bits_active_vidiv & (_T_137 | _T_9);	// sequencer-master.scala:232:25
      wire _T_1781 = io_op_bits_active_vidiv & (_T_138 | _T_10);	// sequencer-master.scala:232:25
      wire _T_1782 = io_op_bits_active_vidiv & (&_T_0 | &tail);	// sequencer-master.scala:232:25, :267:35, util.scala:94:11
      wire [1:0] _io_op_bits_fn_union_7to6 = io_op_bits_fn_union[7:6];	// types-vxu.scala:95:47
      wire _T_1783 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1784 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & _T_1759) : _T_1759;	// sequencer-master.scala:273:29, :329:29
      wire _T_1785 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1786 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1787 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1788 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1789 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & _T_1760) : _T_1760;	// sequencer-master.scala:273:29, :329:29
      wire _T_1790 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1791 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1792 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1793 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1794 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & _T_1761) : _T_1761;	// sequencer-master.scala:273:29, :329:29
      wire _T_1795 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1796 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1797 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1798 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1799 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & _T_1762) : _T_1762;	// sequencer-master.scala:273:29, :329:29
      wire _T_1800 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1801 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1802 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1803 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1804 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & _T_1763) : _T_1763;	// sequencer-master.scala:273:29, :329:29
      wire _T_1805 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1806 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1807 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1808 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1809 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & _T_1764) : _T_1764;	// sequencer-master.scala:273:29, :329:29
      wire _T_1810 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1811 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1812 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1813 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1814 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid :
                ~_T_10 & _T_1765) : _T_1765;	// sequencer-master.scala:273:29, :329:29
      wire _T_1815 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1816 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1817 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1818 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1819 = io_op_bits_active_vfma ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid :
                ~(&tail) & _T_1766) : _T_1766;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1820 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1821 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1822 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1823 = io_op_bits_active_vfma & _T_4;	// sequencer-master.scala:230:21
      wire _T_1824 = io_op_bits_active_vfma & _T_5;	// sequencer-master.scala:230:21
      wire _T_1825 = io_op_bits_active_vfma & _T_6;	// sequencer-master.scala:230:21
      wire _T_1826 = io_op_bits_active_vfma & _T_7;	// sequencer-master.scala:230:21
      wire _T_1827 = io_op_bits_active_vfma & _T_8;	// sequencer-master.scala:230:21
      wire _T_1828 = io_op_bits_active_vfma & _T_9;	// sequencer-master.scala:230:21
      wire _T_1829 = io_op_bits_active_vfma & _T_10;	// sequencer-master.scala:230:21
      wire _T_1830 = io_op_bits_active_vfma & &tail;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [7:0] _T_1831 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1783 ?
                io_op_bits_base_vs1_id : _T_1727) : _T_1783 ? io_op_bits_base_vs1_id : _T_1727;	// sequencer-master.scala:329:29
      wire _T_1832 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1785 ?
                io_op_bits_base_vs1_scalar : _T_1728) : _T_1785 ? io_op_bits_base_vs1_scalar : _T_1728;	// sequencer-master.scala:329:29
      wire _T_1833 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1786 ?
                io_op_bits_base_vs1_pred : _T_1729) : _T_1786 ? io_op_bits_base_vs1_pred : _T_1729;	// sequencer-master.scala:329:29
      wire [1:0] _T_1834 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1787 ?
                io_op_bits_base_vs1_prec : _T_1730) : _T_1787 ? io_op_bits_base_vs1_prec : _T_1730;	// sequencer-master.scala:329:29
      wire [7:0] _T_1835 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1788 ?
                io_op_bits_base_vs1_id : _T_1731) : _T_1788 ? io_op_bits_base_vs1_id : _T_1731;	// sequencer-master.scala:329:29
      wire _T_1836 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1790 ?
                io_op_bits_base_vs1_scalar : _T_1732) : _T_1790 ? io_op_bits_base_vs1_scalar : _T_1732;	// sequencer-master.scala:329:29
      wire _T_1837 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1791 ?
                io_op_bits_base_vs1_pred : _T_1733) : _T_1791 ? io_op_bits_base_vs1_pred : _T_1733;	// sequencer-master.scala:329:29
      wire [1:0] _T_1838 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1792 ?
                io_op_bits_base_vs1_prec : _T_1734) : _T_1792 ? io_op_bits_base_vs1_prec : _T_1734;	// sequencer-master.scala:329:29
      wire [7:0] _T_1839 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1793 ?
                io_op_bits_base_vs1_id : _T_1735) : _T_1793 ? io_op_bits_base_vs1_id : _T_1735;	// sequencer-master.scala:329:29
      wire _T_1840 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1795 ?
                io_op_bits_base_vs1_scalar : _T_1736) : _T_1795 ? io_op_bits_base_vs1_scalar : _T_1736;	// sequencer-master.scala:329:29
      wire _T_1841 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1796 ?
                io_op_bits_base_vs1_pred : _T_1737) : _T_1796 ? io_op_bits_base_vs1_pred : _T_1737;	// sequencer-master.scala:329:29
      wire [1:0] _T_1842 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1797 ?
                io_op_bits_base_vs1_prec : _T_1738) : _T_1797 ? io_op_bits_base_vs1_prec : _T_1738;	// sequencer-master.scala:329:29
      wire [7:0] _T_1843 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1798 ?
                io_op_bits_base_vs1_id : _T_1739) : _T_1798 ? io_op_bits_base_vs1_id : _T_1739;	// sequencer-master.scala:329:29
      wire _T_1844 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1800 ?
                io_op_bits_base_vs1_scalar : _T_1740) : _T_1800 ? io_op_bits_base_vs1_scalar : _T_1740;	// sequencer-master.scala:329:29
      wire _T_1845 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1801 ?
                io_op_bits_base_vs1_pred : _T_1741) : _T_1801 ? io_op_bits_base_vs1_pred : _T_1741;	// sequencer-master.scala:329:29
      wire [1:0] _T_1846 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1802 ?
                io_op_bits_base_vs1_prec : _T_1742) : _T_1802 ? io_op_bits_base_vs1_prec : _T_1742;	// sequencer-master.scala:329:29
      wire [7:0] _T_1847 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1803 ?
                io_op_bits_base_vs1_id : _T_1743) : _T_1803 ? io_op_bits_base_vs1_id : _T_1743;	// sequencer-master.scala:329:29
      wire _T_1848 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1805 ?
                io_op_bits_base_vs1_scalar : _T_1744) : _T_1805 ? io_op_bits_base_vs1_scalar : _T_1744;	// sequencer-master.scala:329:29
      wire _T_1849 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1806 ?
                io_op_bits_base_vs1_pred : _T_1745) : _T_1806 ? io_op_bits_base_vs1_pred : _T_1745;	// sequencer-master.scala:329:29
      wire [1:0] _T_1850 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1807 ?
                io_op_bits_base_vs1_prec : _T_1746) : _T_1807 ? io_op_bits_base_vs1_prec : _T_1746;	// sequencer-master.scala:329:29
      wire [7:0] _T_1851 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1808 ?
                io_op_bits_base_vs1_id : _T_1747) : _T_1808 ? io_op_bits_base_vs1_id : _T_1747;	// sequencer-master.scala:329:29
      wire _T_1852 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1810 ?
                io_op_bits_base_vs1_scalar : _T_1748) : _T_1810 ? io_op_bits_base_vs1_scalar : _T_1748;	// sequencer-master.scala:329:29
      wire _T_1853 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1811 ?
                io_op_bits_base_vs1_pred : _T_1749) : _T_1811 ? io_op_bits_base_vs1_pred : _T_1749;	// sequencer-master.scala:329:29
      wire [1:0] _T_1854 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1812 ?
                io_op_bits_base_vs1_prec : _T_1750) : _T_1812 ? io_op_bits_base_vs1_prec : _T_1750;	// sequencer-master.scala:329:29
      wire [7:0] _T_1855 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1813 ?
                io_op_bits_base_vs1_id : _T_1751) : _T_1813 ? io_op_bits_base_vs1_id : _T_1751;	// sequencer-master.scala:329:29
      wire _T_1856 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1815 ?
                io_op_bits_base_vs1_scalar : _T_1752) : _T_1815 ? io_op_bits_base_vs1_scalar : _T_1752;	// sequencer-master.scala:329:29
      wire _T_1857 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1816 ?
                io_op_bits_base_vs1_pred : _T_1753) : _T_1816 ? io_op_bits_base_vs1_pred : _T_1753;	// sequencer-master.scala:329:29
      wire [1:0] _T_1858 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1817 ?
                io_op_bits_base_vs1_prec : _T_1754) : _T_1817 ? io_op_bits_base_vs1_prec : _T_1754;	// sequencer-master.scala:329:29
      wire [7:0] _T_1859 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (&tail | _T_1818 ?
                io_op_bits_base_vs1_id : _T_1755) : _T_1818 ? io_op_bits_base_vs1_id : _T_1755;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1860 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (&tail | _T_1820 ?
                io_op_bits_base_vs1_scalar : _T_1756) : _T_1820 ? io_op_bits_base_vs1_scalar : _T_1756;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1861 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (&tail | _T_1821 ?
                io_op_bits_base_vs1_pred : _T_1757) : _T_1821 ? io_op_bits_base_vs1_pred : _T_1757;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_1862 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid ? (&tail | _T_1822 ?
                io_op_bits_base_vs1_prec : _T_1758) : _T_1822 ? io_op_bits_base_vs1_prec : _T_1758;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1863 = io_op_bits_active_vfdiv ? ~_T_132 & (io_op_bits_base_vs1_valid & _T_4 ?
                io_op_bits_base_vs1_valid : ~_T_4 & _T_1784) : _T_1784;	// sequencer-master.scala:273:29, :329:29
      wire _T_1864 = io_op_bits_active_vfdiv ? ~_T_133 & (io_op_bits_base_vs1_valid & _T_5 ?
                io_op_bits_base_vs1_valid : ~_T_5 & _T_1789) : _T_1789;	// sequencer-master.scala:273:29, :329:29
      wire _T_1865 = io_op_bits_active_vfdiv ? ~_T_134 & (io_op_bits_base_vs1_valid & _T_6 ?
                io_op_bits_base_vs1_valid : ~_T_6 & _T_1794) : _T_1794;	// sequencer-master.scala:273:29, :329:29
      wire _T_1866 = io_op_bits_active_vfdiv ? ~_T_135 & (io_op_bits_base_vs1_valid & _T_7 ?
                io_op_bits_base_vs1_valid : ~_T_7 & _T_1799) : _T_1799;	// sequencer-master.scala:273:29, :329:29
      wire _T_1867 = io_op_bits_active_vfdiv ? ~_T_136 & (io_op_bits_base_vs1_valid & _T_8 ?
                io_op_bits_base_vs1_valid : ~_T_8 & _T_1804) : _T_1804;	// sequencer-master.scala:273:29, :329:29
      wire _T_1868 = io_op_bits_active_vfdiv ? ~_T_137 & (io_op_bits_base_vs1_valid & _T_9 ?
                io_op_bits_base_vs1_valid : ~_T_9 & _T_1809) : _T_1809;	// sequencer-master.scala:273:29, :329:29
      wire _T_1869 = io_op_bits_active_vfdiv ? ~_T_138 & (io_op_bits_base_vs1_valid & _T_10 ?
                io_op_bits_base_vs1_valid : ~_T_10 & _T_1814) : _T_1814;	// sequencer-master.scala:273:29, :329:29
      wire _T_1870 = io_op_bits_active_vfdiv ? ~(&_T_0) & (io_op_bits_base_vs1_valid & &tail ?
                io_op_bits_base_vs1_valid : ~(&tail) & _T_1819) : _T_1819;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1871 = io_op_bits_active_vfdiv & (_T_132 | _T_4);	// sequencer-master.scala:231:25
      wire _T_1872 = io_op_bits_active_vfdiv & (_T_133 | _T_5);	// sequencer-master.scala:231:25
      wire _T_1873 = io_op_bits_active_vfdiv & (_T_134 | _T_6);	// sequencer-master.scala:231:25
      wire _T_1874 = io_op_bits_active_vfdiv & (_T_135 | _T_7);	// sequencer-master.scala:231:25
      wire _T_1875 = io_op_bits_active_vfdiv & (_T_136 | _T_8);	// sequencer-master.scala:231:25
      wire _T_1876 = io_op_bits_active_vfdiv & (_T_137 | _T_9);	// sequencer-master.scala:231:25
      wire _T_1877 = io_op_bits_active_vfdiv & (_T_138 | _T_10);	// sequencer-master.scala:231:25
      wire _T_1878 = io_op_bits_active_vfdiv & (&_T_0 | &tail);	// sequencer-master.scala:231:25, :267:35, util.scala:94:11
      wire _T_1879 = io_op_bits_active_vfdiv & (_T_132 | _T_4);	// sequencer-master.scala:232:25
      wire _T_1880 = io_op_bits_active_vfdiv & (_T_133 | _T_5);	// sequencer-master.scala:232:25
      wire _T_1881 = io_op_bits_active_vfdiv & (_T_134 | _T_6);	// sequencer-master.scala:232:25
      wire _T_1882 = io_op_bits_active_vfdiv & (_T_135 | _T_7);	// sequencer-master.scala:232:25
      wire _T_1883 = io_op_bits_active_vfdiv & (_T_136 | _T_8);	// sequencer-master.scala:232:25
      wire _T_1884 = io_op_bits_active_vfdiv & (_T_137 | _T_9);	// sequencer-master.scala:232:25
      wire _T_1885 = io_op_bits_active_vfdiv & (_T_138 | _T_10);	// sequencer-master.scala:232:25
      wire _T_1886 = io_op_bits_active_vfdiv & (&_T_0 | &tail);	// sequencer-master.scala:232:25, :267:35, util.scala:94:11
      wire _T_1887 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1888 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & _T_1863) : _T_1863;	// sequencer-master.scala:273:29, :329:29
      wire _T_1889 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1890 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1891 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_1892 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1893 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & _T_1864) : _T_1864;	// sequencer-master.scala:273:29, :329:29
      wire _T_1894 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1895 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1896 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_1897 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1898 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & _T_1865) : _T_1865;	// sequencer-master.scala:273:29, :329:29
      wire _T_1899 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1900 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1901 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_1902 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1903 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & _T_1866) : _T_1866;	// sequencer-master.scala:273:29, :329:29
      wire _T_1904 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1905 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1906 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_1907 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1908 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & _T_1867) : _T_1867;	// sequencer-master.scala:273:29, :329:29
      wire _T_1909 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1910 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1911 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_1912 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1913 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & _T_1868) : _T_1868;	// sequencer-master.scala:273:29, :329:29
      wire _T_1914 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1915 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1916 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_1917 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1918 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid :
                ~_T_10 & _T_1869) : _T_1869;	// sequencer-master.scala:273:29, :329:29
      wire _T_1919 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1920 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1921 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_1922 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1923 = io_op_bits_active_vfcmp ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid :
                ~(&tail) & _T_1870) : _T_1870;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1924 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1925 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1926 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1927 = io_op_bits_active_vfcmp & _T_4;	// sequencer-master.scala:230:21
      wire _T_1928 = io_op_bits_active_vfcmp & _T_5;	// sequencer-master.scala:230:21
      wire _T_1929 = io_op_bits_active_vfcmp & _T_6;	// sequencer-master.scala:230:21
      wire _T_1930 = io_op_bits_active_vfcmp & _T_7;	// sequencer-master.scala:230:21
      wire _T_1931 = io_op_bits_active_vfcmp & _T_8;	// sequencer-master.scala:230:21
      wire _T_1932 = io_op_bits_active_vfcmp & _T_9;	// sequencer-master.scala:230:21
      wire _T_1933 = io_op_bits_active_vfcmp & _T_10;	// sequencer-master.scala:230:21
      wire _T_1934 = io_op_bits_active_vfcmp & &tail;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [7:0] _T_1935 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1887 ?
                io_op_bits_base_vs1_id : _T_1831) : _T_1887 ? io_op_bits_base_vs1_id : _T_1831;	// sequencer-master.scala:329:29
      wire _T_1936 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1889 ?
                io_op_bits_base_vs1_scalar : _T_1832) : _T_1889 ? io_op_bits_base_vs1_scalar : _T_1832;	// sequencer-master.scala:329:29
      wire _T_1937 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1890 ?
                io_op_bits_base_vs1_pred : _T_1833) : _T_1890 ? io_op_bits_base_vs1_pred : _T_1833;	// sequencer-master.scala:329:29
      wire [1:0] _T_1938 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_4 | _T_1891 ?
                io_op_bits_base_vs1_prec : _T_1834) : _T_1891 ? io_op_bits_base_vs1_prec : _T_1834;	// sequencer-master.scala:329:29
      wire [7:0] _T_1939 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1892 ?
                io_op_bits_base_vs1_id : _T_1835) : _T_1892 ? io_op_bits_base_vs1_id : _T_1835;	// sequencer-master.scala:329:29
      wire _T_1940 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1894 ?
                io_op_bits_base_vs1_scalar : _T_1836) : _T_1894 ? io_op_bits_base_vs1_scalar : _T_1836;	// sequencer-master.scala:329:29
      wire _T_1941 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1895 ?
                io_op_bits_base_vs1_pred : _T_1837) : _T_1895 ? io_op_bits_base_vs1_pred : _T_1837;	// sequencer-master.scala:329:29
      wire [1:0] _T_1942 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_5 | _T_1896 ?
                io_op_bits_base_vs1_prec : _T_1838) : _T_1896 ? io_op_bits_base_vs1_prec : _T_1838;	// sequencer-master.scala:329:29
      wire [7:0] _T_1943 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1897 ?
                io_op_bits_base_vs1_id : _T_1839) : _T_1897 ? io_op_bits_base_vs1_id : _T_1839;	// sequencer-master.scala:329:29
      wire _T_1944 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1899 ?
                io_op_bits_base_vs1_scalar : _T_1840) : _T_1899 ? io_op_bits_base_vs1_scalar : _T_1840;	// sequencer-master.scala:329:29
      wire _T_1945 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1900 ?
                io_op_bits_base_vs1_pred : _T_1841) : _T_1900 ? io_op_bits_base_vs1_pred : _T_1841;	// sequencer-master.scala:329:29
      wire [1:0] _T_1946 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_6 | _T_1901 ?
                io_op_bits_base_vs1_prec : _T_1842) : _T_1901 ? io_op_bits_base_vs1_prec : _T_1842;	// sequencer-master.scala:329:29
      wire [7:0] _T_1947 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1902 ?
                io_op_bits_base_vs1_id : _T_1843) : _T_1902 ? io_op_bits_base_vs1_id : _T_1843;	// sequencer-master.scala:329:29
      wire _T_1948 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1904 ?
                io_op_bits_base_vs1_scalar : _T_1844) : _T_1904 ? io_op_bits_base_vs1_scalar : _T_1844;	// sequencer-master.scala:329:29
      wire _T_1949 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1905 ?
                io_op_bits_base_vs1_pred : _T_1845) : _T_1905 ? io_op_bits_base_vs1_pred : _T_1845;	// sequencer-master.scala:329:29
      wire [1:0] _T_1950 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_7 | _T_1906 ?
                io_op_bits_base_vs1_prec : _T_1846) : _T_1906 ? io_op_bits_base_vs1_prec : _T_1846;	// sequencer-master.scala:329:29
      wire [7:0] _T_1951 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1907 ?
                io_op_bits_base_vs1_id : _T_1847) : _T_1907 ? io_op_bits_base_vs1_id : _T_1847;	// sequencer-master.scala:329:29
      wire _T_1952 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1909 ?
                io_op_bits_base_vs1_scalar : _T_1848) : _T_1909 ? io_op_bits_base_vs1_scalar : _T_1848;	// sequencer-master.scala:329:29
      wire _T_1953 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1910 ?
                io_op_bits_base_vs1_pred : _T_1849) : _T_1910 ? io_op_bits_base_vs1_pred : _T_1849;	// sequencer-master.scala:329:29
      wire [1:0] _T_1954 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_8 | _T_1911 ?
                io_op_bits_base_vs1_prec : _T_1850) : _T_1911 ? io_op_bits_base_vs1_prec : _T_1850;	// sequencer-master.scala:329:29
      wire [7:0] _T_1955 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1912 ?
                io_op_bits_base_vs1_id : _T_1851) : _T_1912 ? io_op_bits_base_vs1_id : _T_1851;	// sequencer-master.scala:329:29
      wire _T_1956 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1914 ?
                io_op_bits_base_vs1_scalar : _T_1852) : _T_1914 ? io_op_bits_base_vs1_scalar : _T_1852;	// sequencer-master.scala:329:29
      wire _T_1957 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1915 ?
                io_op_bits_base_vs1_pred : _T_1853) : _T_1915 ? io_op_bits_base_vs1_pred : _T_1853;	// sequencer-master.scala:329:29
      wire [1:0] _T_1958 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_9 | _T_1916 ?
                io_op_bits_base_vs1_prec : _T_1854) : _T_1916 ? io_op_bits_base_vs1_prec : _T_1854;	// sequencer-master.scala:329:29
      wire [7:0] _T_1959 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1917 ?
                io_op_bits_base_vs1_id : _T_1855) : _T_1917 ? io_op_bits_base_vs1_id : _T_1855;	// sequencer-master.scala:329:29
      wire _T_1960 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1919 ?
                io_op_bits_base_vs1_scalar : _T_1856) : _T_1919 ? io_op_bits_base_vs1_scalar : _T_1856;	// sequencer-master.scala:329:29
      wire _T_1961 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1920 ?
                io_op_bits_base_vs1_pred : _T_1857) : _T_1920 ? io_op_bits_base_vs1_pred : _T_1857;	// sequencer-master.scala:329:29
      wire [1:0] _T_1962 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (_T_10 | _T_1921 ?
                io_op_bits_base_vs1_prec : _T_1858) : _T_1921 ? io_op_bits_base_vs1_prec : _T_1858;	// sequencer-master.scala:329:29
      wire [7:0] _T_1963 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (&tail | _T_1922 ?
                io_op_bits_base_vs1_id : _T_1859) : _T_1922 ? io_op_bits_base_vs1_id : _T_1859;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1964 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (&tail | _T_1924 ?
                io_op_bits_base_vs1_scalar : _T_1860) : _T_1924 ? io_op_bits_base_vs1_scalar : _T_1860;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1965 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (&tail | _T_1925 ?
                io_op_bits_base_vs1_pred : _T_1861) : _T_1925 ? io_op_bits_base_vs1_pred : _T_1861;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_1966 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid ? (&tail | _T_1926 ?
                io_op_bits_base_vs1_prec : _T_1862) : _T_1926 ? io_op_bits_base_vs1_prec : _T_1862;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_1967 = (~io_op_bits_active_vrpred | ~_T_4) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid : ~_T_4 & _T_1888) : _T_1888);	// sequencer-master.scala:273:29, :329:29
      wire _T_1968 = (~io_op_bits_active_vrpred | ~_T_5) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid : ~_T_5 & _T_1893) : _T_1893);	// sequencer-master.scala:273:29, :329:29
      wire _T_1969 = (~io_op_bits_active_vrpred | ~_T_6) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid : ~_T_6 & _T_1898) : _T_1898);	// sequencer-master.scala:273:29, :329:29
      wire _T_1970 = (~io_op_bits_active_vrpred | ~_T_7) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid : ~_T_7 & _T_1903) : _T_1903);	// sequencer-master.scala:273:29, :329:29
      wire _T_1971 = (~io_op_bits_active_vrpred | ~_T_8) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid : ~_T_8 & _T_1908) : _T_1908);	// sequencer-master.scala:273:29, :329:29
      wire _T_1972 = (~io_op_bits_active_vrpred | ~_T_9) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid : ~_T_9 & _T_1913) : _T_1913);	// sequencer-master.scala:273:29, :329:29
      wire _T_1973 = (~io_op_bits_active_vrpred | ~_T_10) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid : ~_T_10 & _T_1918) :
                _T_1918);	// sequencer-master.scala:273:29, :329:29
      wire _T_1974 = (~io_op_bits_active_vrpred | ~(&tail)) & (io_op_bits_active_vfconv ?
                (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid : ~(&tail) & _T_1923) :
                _T_1923);	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_1975 = io_op_bits_active_vrpred & _T_4;	// sequencer-master.scala:230:21
      wire _T_1976 = io_op_bits_active_vrpred & _T_5;	// sequencer-master.scala:230:21
      wire _T_1977 = io_op_bits_active_vrpred & _T_6;	// sequencer-master.scala:230:21
      wire _T_1978 = io_op_bits_active_vrpred & _T_7;	// sequencer-master.scala:230:21
      wire _T_1979 = io_op_bits_active_vrpred & _T_8;	// sequencer-master.scala:230:21
      wire _T_1980 = io_op_bits_active_vrpred & _T_9;	// sequencer-master.scala:230:21
      wire _T_1981 = io_op_bits_active_vrpred & _T_10;	// sequencer-master.scala:230:21
      wire _T_1982 = io_op_bits_active_vrpred & &tail;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire _T_1983 = io_op_bits_active_vrpred & _T_4;	// sequencer-master.scala:231:25
      wire _T_1984 = io_op_bits_active_vrpred & _T_5;	// sequencer-master.scala:231:25
      wire _T_1985 = io_op_bits_active_vrpred & _T_6;	// sequencer-master.scala:231:25
      wire _T_1986 = io_op_bits_active_vrpred & _T_7;	// sequencer-master.scala:231:25
      wire _T_1987 = io_op_bits_active_vrpred & _T_8;	// sequencer-master.scala:231:25
      wire _T_1988 = io_op_bits_active_vrpred & _T_9;	// sequencer-master.scala:231:25
      wire _T_1989 = io_op_bits_active_vrpred & _T_10;	// sequencer-master.scala:231:25
      wire _T_1990 = io_op_bits_active_vrpred & &tail;	// sequencer-master.scala:231:25, :267:35, util.scala:94:11
      wire _T_1991 = io_op_bits_active_vrpred & _T_4;	// sequencer-master.scala:232:25
      wire _T_1992 = io_op_bits_active_vrpred & _T_5;	// sequencer-master.scala:232:25
      wire _T_1993 = io_op_bits_active_vrpred & _T_6;	// sequencer-master.scala:232:25
      wire _T_1994 = io_op_bits_active_vrpred & _T_7;	// sequencer-master.scala:232:25
      wire _T_1995 = io_op_bits_active_vrpred & _T_8;	// sequencer-master.scala:232:25
      wire _T_1996 = io_op_bits_active_vrpred & _T_9;	// sequencer-master.scala:232:25
      wire _T_1997 = io_op_bits_active_vrpred & _T_10;	// sequencer-master.scala:232:25
      wire _T_1998 = io_op_bits_active_vrpred & &tail;	// sequencer-master.scala:232:25, :267:35, util.scala:94:11
      wire _T_1999 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire [7:0] _T_2000 = _T_1999 ? io_op_bits_base_vs1_id : _T_1935;	// sequencer-master.scala:329:29
      wire _T_2001 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_4 ? io_op_bits_base_vs1_valid :
                ~_T_4 & _T_1967) : _T_1967;	// sequencer-master.scala:273:29, :329:29
      wire _T_2002 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_2003 = _T_2002 ? io_op_bits_base_vs1_scalar : _T_1936;	// sequencer-master.scala:329:29
      wire _T_2004 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_2005 = _T_2004 ? io_op_bits_base_vs1_pred : _T_1937;	// sequencer-master.scala:329:29
      wire _T_2006 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_4;	// sequencer-master.scala:329:29
      wire [1:0] _T_2007 = _T_2006 ? io_op_bits_base_vs1_prec : _T_1938;	// sequencer-master.scala:329:29
      wire _T_2008 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire [7:0] _T_2009 = _T_2008 ? io_op_bits_base_vs1_id : _T_1939;	// sequencer-master.scala:329:29
      wire _T_2010 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_5 ? io_op_bits_base_vs1_valid :
                ~_T_5 & _T_1968) : _T_1968;	// sequencer-master.scala:273:29, :329:29
      wire _T_2011 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_2012 = _T_2011 ? io_op_bits_base_vs1_scalar : _T_1940;	// sequencer-master.scala:329:29
      wire _T_2013 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_2014 = _T_2013 ? io_op_bits_base_vs1_pred : _T_1941;	// sequencer-master.scala:329:29
      wire _T_2015 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_5;	// sequencer-master.scala:329:29
      wire [1:0] _T_2016 = _T_2015 ? io_op_bits_base_vs1_prec : _T_1942;	// sequencer-master.scala:329:29
      wire _T_2017 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire [7:0] _T_2018 = _T_2017 ? io_op_bits_base_vs1_id : _T_1943;	// sequencer-master.scala:329:29
      wire _T_2019 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_6 ? io_op_bits_base_vs1_valid :
                ~_T_6 & _T_1969) : _T_1969;	// sequencer-master.scala:273:29, :329:29
      wire _T_2020 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_2021 = _T_2020 ? io_op_bits_base_vs1_scalar : _T_1944;	// sequencer-master.scala:329:29
      wire _T_2022 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_2023 = _T_2022 ? io_op_bits_base_vs1_pred : _T_1945;	// sequencer-master.scala:329:29
      wire _T_2024 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_6;	// sequencer-master.scala:329:29
      wire [1:0] _T_2025 = _T_2024 ? io_op_bits_base_vs1_prec : _T_1946;	// sequencer-master.scala:329:29
      wire _T_2026 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire [7:0] _T_2027 = _T_2026 ? io_op_bits_base_vs1_id : _T_1947;	// sequencer-master.scala:329:29
      wire _T_2028 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_7 ? io_op_bits_base_vs1_valid :
                ~_T_7 & _T_1970) : _T_1970;	// sequencer-master.scala:273:29, :329:29
      wire _T_2029 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_2030 = _T_2029 ? io_op_bits_base_vs1_scalar : _T_1948;	// sequencer-master.scala:329:29
      wire _T_2031 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_2032 = _T_2031 ? io_op_bits_base_vs1_pred : _T_1949;	// sequencer-master.scala:329:29
      wire _T_2033 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_7;	// sequencer-master.scala:329:29
      wire [1:0] _T_2034 = _T_2033 ? io_op_bits_base_vs1_prec : _T_1950;	// sequencer-master.scala:329:29
      wire _T_2035 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire [7:0] _T_2036 = _T_2035 ? io_op_bits_base_vs1_id : _T_1951;	// sequencer-master.scala:329:29
      wire _T_2037 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_8 ? io_op_bits_base_vs1_valid :
                ~_T_8 & _T_1971) : _T_1971;	// sequencer-master.scala:273:29, :329:29
      wire _T_2038 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_2039 = _T_2038 ? io_op_bits_base_vs1_scalar : _T_1952;	// sequencer-master.scala:329:29
      wire _T_2040 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_2041 = _T_2040 ? io_op_bits_base_vs1_pred : _T_1953;	// sequencer-master.scala:329:29
      wire _T_2042 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_8;	// sequencer-master.scala:329:29
      wire [1:0] _T_2043 = _T_2042 ? io_op_bits_base_vs1_prec : _T_1954;	// sequencer-master.scala:329:29
      wire _T_2044 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire [7:0] _T_2045 = _T_2044 ? io_op_bits_base_vs1_id : _T_1955;	// sequencer-master.scala:329:29
      wire _T_2046 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_9 ? io_op_bits_base_vs1_valid :
                ~_T_9 & _T_1972) : _T_1972;	// sequencer-master.scala:273:29, :329:29
      wire _T_2047 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_2048 = _T_2047 ? io_op_bits_base_vs1_scalar : _T_1956;	// sequencer-master.scala:329:29
      wire _T_2049 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_2050 = _T_2049 ? io_op_bits_base_vs1_pred : _T_1957;	// sequencer-master.scala:329:29
      wire _T_2051 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_9;	// sequencer-master.scala:329:29
      wire [1:0] _T_2052 = _T_2051 ? io_op_bits_base_vs1_prec : _T_1958;	// sequencer-master.scala:329:29
      wire _T_2053 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire [7:0] _T_2054 = _T_2053 ? io_op_bits_base_vs1_id : _T_1959;	// sequencer-master.scala:329:29
      wire _T_2055 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & _T_10 ? io_op_bits_base_vs1_valid
                : ~_T_10 & _T_1973) : _T_1973;	// sequencer-master.scala:273:29, :329:29
      wire _T_2056 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_2057 = _T_2056 ? io_op_bits_base_vs1_scalar : _T_1960;	// sequencer-master.scala:329:29
      wire _T_2058 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_2059 = _T_2058 ? io_op_bits_base_vs1_pred : _T_1961;	// sequencer-master.scala:329:29
      wire _T_2060 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_10;	// sequencer-master.scala:329:29
      wire [1:0] _T_2061 = _T_2060 ? io_op_bits_base_vs1_prec : _T_1962;	// sequencer-master.scala:329:29
      wire _T_2062 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [7:0] _T_2063 = _T_2062 ? io_op_bits_base_vs1_id : _T_1963;	// sequencer-master.scala:329:29
      wire _T_2064 = io_op_bits_active_vrfirst ? (io_op_bits_base_vs1_valid & &tail ? io_op_bits_base_vs1_valid
                : ~(&tail) & _T_1974) : _T_1974;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_2065 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2066 = _T_2065 ? io_op_bits_base_vs1_scalar : _T_1964;	// sequencer-master.scala:329:29
      wire _T_2067 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2068 = _T_2067 ? io_op_bits_base_vs1_pred : _T_1965;	// sequencer-master.scala:329:29
      wire _T_2069 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_2070 = _T_2069 ? io_op_bits_base_vs1_prec : _T_1966;	// sequencer-master.scala:329:29
      wire [7:0] _T_2071 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_291 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_4 | _T_1999 ? io_op_bits_base_vs1_id : _T_1935) : _T_2000)
                : _T_2000;	// sequencer-master.scala:329:29
      wire _T_2072 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_291 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_4 | _T_2002 ? io_op_bits_base_vs1_scalar : _T_1936) :
                _T_2003) : _T_2003;	// sequencer-master.scala:329:29
      wire _T_2073 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_291 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_4 | _T_2004 ? io_op_bits_base_vs1_pred : _T_1937) :
                _T_2005) : _T_2005;	// sequencer-master.scala:329:29
      wire [1:0] _T_2074 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_291 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_4 | _T_2006 ? io_op_bits_base_vs1_prec : _T_1938) :
                _T_2007) : _T_2007;	// sequencer-master.scala:329:29
      wire [7:0] _T_2075 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_292 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_5 | _T_2008 ? io_op_bits_base_vs1_id : _T_1939) : _T_2009)
                : _T_2009;	// sequencer-master.scala:329:29
      wire _T_2076 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_292 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_5 | _T_2011 ? io_op_bits_base_vs1_scalar : _T_1940) :
                _T_2012) : _T_2012;	// sequencer-master.scala:329:29
      wire _T_2077 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_292 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_5 | _T_2013 ? io_op_bits_base_vs1_pred : _T_1941) :
                _T_2014) : _T_2014;	// sequencer-master.scala:329:29
      wire [1:0] _T_2078 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_292 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_5 | _T_2015 ? io_op_bits_base_vs1_prec : _T_1942) :
                _T_2016) : _T_2016;	// sequencer-master.scala:329:29
      wire [7:0] _T_2079 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_293 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_6 | _T_2017 ? io_op_bits_base_vs1_id : _T_1943) : _T_2018)
                : _T_2018;	// sequencer-master.scala:329:29
      wire _T_2080 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_293 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_6 | _T_2020 ? io_op_bits_base_vs1_scalar : _T_1944) :
                _T_2021) : _T_2021;	// sequencer-master.scala:329:29
      wire _T_2081 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_293 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_6 | _T_2022 ? io_op_bits_base_vs1_pred : _T_1945) :
                _T_2023) : _T_2023;	// sequencer-master.scala:329:29
      wire [1:0] _T_2082 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_293 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_6 | _T_2024 ? io_op_bits_base_vs1_prec : _T_1946) :
                _T_2025) : _T_2025;	// sequencer-master.scala:329:29
      wire [7:0] _T_2083 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_294 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_7 | _T_2026 ? io_op_bits_base_vs1_id : _T_1947) : _T_2027)
                : _T_2027;	// sequencer-master.scala:329:29
      wire _T_2084 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_294 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_7 | _T_2029 ? io_op_bits_base_vs1_scalar : _T_1948) :
                _T_2030) : _T_2030;	// sequencer-master.scala:329:29
      wire _T_2085 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_294 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_7 | _T_2031 ? io_op_bits_base_vs1_pred : _T_1949) :
                _T_2032) : _T_2032;	// sequencer-master.scala:329:29
      wire [1:0] _T_2086 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_294 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_7 | _T_2033 ? io_op_bits_base_vs1_prec : _T_1950) :
                _T_2034) : _T_2034;	// sequencer-master.scala:329:29
      wire [7:0] _T_2087 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_295 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_8 | _T_2035 ? io_op_bits_base_vs1_id : _T_1951) : _T_2036)
                : _T_2036;	// sequencer-master.scala:329:29
      wire _T_2088 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_295 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_8 | _T_2038 ? io_op_bits_base_vs1_scalar : _T_1952) :
                _T_2039) : _T_2039;	// sequencer-master.scala:329:29
      wire _T_2089 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_295 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_8 | _T_2040 ? io_op_bits_base_vs1_pred : _T_1953) :
                _T_2041) : _T_2041;	// sequencer-master.scala:329:29
      wire [1:0] _T_2090 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_295 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_8 | _T_2042 ? io_op_bits_base_vs1_prec : _T_1954) :
                _T_2043) : _T_2043;	// sequencer-master.scala:329:29
      wire [7:0] _T_2091 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_296 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_9 | _T_2044 ? io_op_bits_base_vs1_id : _T_1955) : _T_2045)
                : _T_2045;	// sequencer-master.scala:329:29
      wire _T_2092 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_296 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_9 | _T_2047 ? io_op_bits_base_vs1_scalar : _T_1956) :
                _T_2048) : _T_2048;	// sequencer-master.scala:329:29
      wire _T_2093 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_296 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_9 | _T_2049 ? io_op_bits_base_vs1_pred : _T_1957) :
                _T_2050) : _T_2050;	// sequencer-master.scala:329:29
      wire [1:0] _T_2094 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_296 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_9 | _T_2051 ? io_op_bits_base_vs1_prec : _T_1958) :
                _T_2052) : _T_2052;	// sequencer-master.scala:329:29
      wire [7:0] _T_2095 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_297 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (_T_10 | _T_2053 ? io_op_bits_base_vs1_id : _T_1959) : _T_2054)
                : _T_2054;	// sequencer-master.scala:329:29
      wire _T_2096 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_297 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (_T_10 | _T_2056 ? io_op_bits_base_vs1_scalar : _T_1960) :
                _T_2057) : _T_2057;	// sequencer-master.scala:329:29
      wire _T_2097 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_297 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (_T_10 | _T_2058 ? io_op_bits_base_vs1_pred : _T_1961) :
                _T_2059) : _T_2059;	// sequencer-master.scala:329:29
      wire [1:0] _T_2098 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_297 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (_T_10 | _T_2060 ? io_op_bits_base_vs1_prec : _T_1962) :
                _T_2061) : _T_2061;	// sequencer-master.scala:329:29
      wire [7:0] _T_2099 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & &_T_1 ? io_op_bits_base_vs2_id :
                io_op_bits_base_vs1_valid ? (&tail | _T_2062 ? io_op_bits_base_vs1_id : _T_1963) : _T_2063)
                : _T_2063;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2100 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & &_T_1 ? io_op_bits_base_vs2_scalar :
                io_op_bits_base_vs1_valid ? (&tail | _T_2065 ? io_op_bits_base_vs1_scalar : _T_1964) :
                _T_2066) : _T_2066;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2101 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & &_T_1 ? io_op_bits_base_vs2_pred :
                io_op_bits_base_vs1_valid ? (&tail | _T_2067 ? io_op_bits_base_vs1_pred : _T_1965) :
                _T_2068) : _T_2068;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_2102 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & &_T_1 ? io_op_bits_base_vs2_prec :
                io_op_bits_base_vs1_valid ? (&tail | _T_2069 ? io_op_bits_base_vs1_prec : _T_1966) :
                _T_2070) : _T_2070;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2103 = io_op_bits_active_vamo ? ~_T_314 & (io_op_bits_base_vs2_valid & _T_291 ?
                io_op_bits_base_vs2_valid : ~_T_291 & ~_T_132 & (io_op_bits_base_vs1_valid & _T_4 ?
                io_op_bits_base_vs1_valid : ~_T_4 & _T_2001)) : _T_2001;	// sequencer-master.scala:273:29, :329:29
      wire _T_2104 = io_op_bits_active_vamo ? ~_T_315 & (io_op_bits_base_vs2_valid & _T_292 ?
                io_op_bits_base_vs2_valid : ~_T_292 & ~_T_133 & (io_op_bits_base_vs1_valid & _T_5 ?
                io_op_bits_base_vs1_valid : ~_T_5 & _T_2010)) : _T_2010;	// sequencer-master.scala:273:29, :329:29
      wire _T_2105 = io_op_bits_active_vamo ? ~_T_316 & (io_op_bits_base_vs2_valid & _T_293 ?
                io_op_bits_base_vs2_valid : ~_T_293 & ~_T_134 & (io_op_bits_base_vs1_valid & _T_6 ?
                io_op_bits_base_vs1_valid : ~_T_6 & _T_2019)) : _T_2019;	// sequencer-master.scala:273:29, :329:29
      wire _T_2106 = io_op_bits_active_vamo ? ~_T_317 & (io_op_bits_base_vs2_valid & _T_294 ?
                io_op_bits_base_vs2_valid : ~_T_294 & ~_T_135 & (io_op_bits_base_vs1_valid & _T_7 ?
                io_op_bits_base_vs1_valid : ~_T_7 & _T_2028)) : _T_2028;	// sequencer-master.scala:273:29, :329:29
      wire _T_2107 = io_op_bits_active_vamo ? ~_T_318 & (io_op_bits_base_vs2_valid & _T_295 ?
                io_op_bits_base_vs2_valid : ~_T_295 & ~_T_136 & (io_op_bits_base_vs1_valid & _T_8 ?
                io_op_bits_base_vs1_valid : ~_T_8 & _T_2037)) : _T_2037;	// sequencer-master.scala:273:29, :329:29
      wire _T_2108 = io_op_bits_active_vamo ? ~_T_319 & (io_op_bits_base_vs2_valid & _T_296 ?
                io_op_bits_base_vs2_valid : ~_T_296 & ~_T_137 & (io_op_bits_base_vs1_valid & _T_9 ?
                io_op_bits_base_vs1_valid : ~_T_9 & _T_2046)) : _T_2046;	// sequencer-master.scala:273:29, :329:29
      wire _T_2109 = io_op_bits_active_vamo ? ~_T_320 & (io_op_bits_base_vs2_valid & _T_297 ?
                io_op_bits_base_vs2_valid : ~_T_297 & ~_T_138 & (io_op_bits_base_vs1_valid & _T_10 ?
                io_op_bits_base_vs1_valid : ~_T_10 & _T_2055)) : _T_2055;	// sequencer-master.scala:273:29, :329:29
      wire _T_2110 = io_op_bits_active_vamo ? ~(&_T_2) & (io_op_bits_base_vs2_valid & &_T_1 ?
                io_op_bits_base_vs2_valid : ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vs1_valid & &tail ?
                io_op_bits_base_vs1_valid : ~(&tail) & _T_2064)) : _T_2064;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_2111 = io_op_bits_active_vamo & (_T_314 | _T_291 | _T_132 | _T_4);	// sequencer-master.scala:231:25
      wire _T_2112 = io_op_bits_active_vamo & (_T_315 | _T_292 | _T_133 | _T_5);	// sequencer-master.scala:231:25
      wire _T_2113 = io_op_bits_active_vamo & (_T_316 | _T_293 | _T_134 | _T_6);	// sequencer-master.scala:231:25
      wire _T_2114 = io_op_bits_active_vamo & (_T_317 | _T_294 | _T_135 | _T_7);	// sequencer-master.scala:231:25
      wire _T_2115 = io_op_bits_active_vamo & (_T_318 | _T_295 | _T_136 | _T_8);	// sequencer-master.scala:231:25
      wire _T_2116 = io_op_bits_active_vamo & (_T_319 | _T_296 | _T_137 | _T_9);	// sequencer-master.scala:231:25
      wire _T_2117 = io_op_bits_active_vamo & (_T_320 | _T_297 | _T_138 | _T_10);	// sequencer-master.scala:231:25
      wire _T_2118 = io_op_bits_active_vamo & (&_T_2 | &_T_1 | &_T_0 | &tail);	// sequencer-master.scala:231:25, :267:35, util.scala:94:11
      wire _T_2119 = io_op_bits_active_vamo & (_T_314 | _T_291 | _T_132 | _T_4);	// sequencer-master.scala:232:25
      wire _T_2120 = io_op_bits_active_vamo & (_T_315 | _T_292 | _T_133 | _T_5);	// sequencer-master.scala:232:25
      wire _T_2121 = io_op_bits_active_vamo & (_T_316 | _T_293 | _T_134 | _T_6);	// sequencer-master.scala:232:25
      wire _T_2122 = io_op_bits_active_vamo & (_T_317 | _T_294 | _T_135 | _T_7);	// sequencer-master.scala:232:25
      wire _T_2123 = io_op_bits_active_vamo & (_T_318 | _T_295 | _T_136 | _T_8);	// sequencer-master.scala:232:25
      wire _T_2124 = io_op_bits_active_vamo & (_T_319 | _T_296 | _T_137 | _T_9);	// sequencer-master.scala:232:25
      wire _T_2125 = io_op_bits_active_vamo & (_T_320 | _T_297 | _T_138 | _T_10);	// sequencer-master.scala:232:25
      wire _T_2126 = io_op_bits_active_vamo & (&_T_2 | &_T_1 | &_T_0 | &tail);	// sequencer-master.scala:232:25, :267:35, util.scala:94:11
      wire _T_2127 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire [7:0] _T_2128 = _T_2127 ? io_op_bits_base_vs2_id : _T_2071;	// sequencer-master.scala:329:29
      wire _T_2129 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_2130 = _T_2129 ? io_op_bits_base_vs2_scalar : _T_2072;	// sequencer-master.scala:329:29
      wire _T_2131 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire _T_2132 = _T_2131 ? io_op_bits_base_vs2_pred : _T_2073;	// sequencer-master.scala:329:29
      wire _T_2133 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_4;	// sequencer-master.scala:329:29
      wire [1:0] _T_2134 = _T_2133 ? io_op_bits_base_vs2_prec : _T_2074;	// sequencer-master.scala:329:29
      wire _T_2135 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire [7:0] _T_2136 = _T_2135 ? io_op_bits_base_vs2_id : _T_2075;	// sequencer-master.scala:329:29
      wire _T_2137 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_2138 = _T_2137 ? io_op_bits_base_vs2_scalar : _T_2076;	// sequencer-master.scala:329:29
      wire _T_2139 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire _T_2140 = _T_2139 ? io_op_bits_base_vs2_pred : _T_2077;	// sequencer-master.scala:329:29
      wire _T_2141 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_5;	// sequencer-master.scala:329:29
      wire [1:0] _T_2142 = _T_2141 ? io_op_bits_base_vs2_prec : _T_2078;	// sequencer-master.scala:329:29
      wire _T_2143 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire [7:0] _T_2144 = _T_2143 ? io_op_bits_base_vs2_id : _T_2079;	// sequencer-master.scala:329:29
      wire _T_2145 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_2146 = _T_2145 ? io_op_bits_base_vs2_scalar : _T_2080;	// sequencer-master.scala:329:29
      wire _T_2147 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire _T_2148 = _T_2147 ? io_op_bits_base_vs2_pred : _T_2081;	// sequencer-master.scala:329:29
      wire _T_2149 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_6;	// sequencer-master.scala:329:29
      wire [1:0] _T_2150 = _T_2149 ? io_op_bits_base_vs2_prec : _T_2082;	// sequencer-master.scala:329:29
      wire _T_2151 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire [7:0] _T_2152 = _T_2151 ? io_op_bits_base_vs2_id : _T_2083;	// sequencer-master.scala:329:29
      wire _T_2153 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_2154 = _T_2153 ? io_op_bits_base_vs2_scalar : _T_2084;	// sequencer-master.scala:329:29
      wire _T_2155 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire _T_2156 = _T_2155 ? io_op_bits_base_vs2_pred : _T_2085;	// sequencer-master.scala:329:29
      wire _T_2157 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_7;	// sequencer-master.scala:329:29
      wire [1:0] _T_2158 = _T_2157 ? io_op_bits_base_vs2_prec : _T_2086;	// sequencer-master.scala:329:29
      wire _T_2159 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire [7:0] _T_2160 = _T_2159 ? io_op_bits_base_vs2_id : _T_2087;	// sequencer-master.scala:329:29
      wire _T_2161 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_2162 = _T_2161 ? io_op_bits_base_vs2_scalar : _T_2088;	// sequencer-master.scala:329:29
      wire _T_2163 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire _T_2164 = _T_2163 ? io_op_bits_base_vs2_pred : _T_2089;	// sequencer-master.scala:329:29
      wire _T_2165 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_8;	// sequencer-master.scala:329:29
      wire [1:0] _T_2166 = _T_2165 ? io_op_bits_base_vs2_prec : _T_2090;	// sequencer-master.scala:329:29
      wire _T_2167 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire [7:0] _T_2168 = _T_2167 ? io_op_bits_base_vs2_id : _T_2091;	// sequencer-master.scala:329:29
      wire _T_2169 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_2170 = _T_2169 ? io_op_bits_base_vs2_scalar : _T_2092;	// sequencer-master.scala:329:29
      wire _T_2171 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire _T_2172 = _T_2171 ? io_op_bits_base_vs2_pred : _T_2093;	// sequencer-master.scala:329:29
      wire _T_2173 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_9;	// sequencer-master.scala:329:29
      wire [1:0] _T_2174 = _T_2173 ? io_op_bits_base_vs2_prec : _T_2094;	// sequencer-master.scala:329:29
      wire _T_2175 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire [7:0] _T_2176 = _T_2175 ? io_op_bits_base_vs2_id : _T_2095;	// sequencer-master.scala:329:29
      wire _T_2177 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_2178 = _T_2177 ? io_op_bits_base_vs2_scalar : _T_2096;	// sequencer-master.scala:329:29
      wire _T_2179 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire _T_2180 = _T_2179 ? io_op_bits_base_vs2_pred : _T_2097;	// sequencer-master.scala:329:29
      wire _T_2181 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_10;	// sequencer-master.scala:329:29
      wire [1:0] _T_2182 = _T_2181 ? io_op_bits_base_vs2_prec : _T_2098;	// sequencer-master.scala:329:29
      wire _T_2183 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [7:0] _T_2184 = _T_2183 ? io_op_bits_base_vs2_id : _T_2099;	// sequencer-master.scala:329:29
      wire _T_2185 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2186 = _T_2185 ? io_op_bits_base_vs2_scalar : _T_2100;	// sequencer-master.scala:329:29
      wire _T_2187 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire _T_2188 = _T_2187 ? io_op_bits_base_vs2_pred : _T_2101;	// sequencer-master.scala:329:29
      wire _T_2189 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & &tail;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      wire [1:0] _T_2190 = _T_2189 ? io_op_bits_base_vs2_prec : _T_2102;	// sequencer-master.scala:329:29
      wire _T_2191 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (io_op_bits_base_vs2_valid & _T_4 ?
                io_op_bits_base_vs2_valid : ~_T_4 & _T_2103) : _T_2103;	// sequencer-master.scala:273:29, :329:29
      wire _T_2192 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (io_op_bits_base_vs2_valid & _T_5 ?
                io_op_bits_base_vs2_valid : ~_T_5 & _T_2104) : _T_2104;	// sequencer-master.scala:273:29, :329:29
      wire _T_2193 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (io_op_bits_base_vs2_valid & _T_6 ?
                io_op_bits_base_vs2_valid : ~_T_6 & _T_2105) : _T_2105;	// sequencer-master.scala:273:29, :329:29
      wire _T_2194 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (io_op_bits_base_vs2_valid & _T_7 ?
                io_op_bits_base_vs2_valid : ~_T_7 & _T_2106) : _T_2106;	// sequencer-master.scala:273:29, :329:29
      wire _T_2195 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (io_op_bits_base_vs2_valid & _T_8 ?
                io_op_bits_base_vs2_valid : ~_T_8 & _T_2107) : _T_2107;	// sequencer-master.scala:273:29, :329:29
      wire _T_2196 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (io_op_bits_base_vs2_valid & _T_9 ?
                io_op_bits_base_vs2_valid : ~_T_9 & _T_2108) : _T_2108;	// sequencer-master.scala:273:29, :329:29
      wire _T_2197 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (io_op_bits_base_vs2_valid & _T_10 ?
                io_op_bits_base_vs2_valid : ~_T_10 & _T_2109) : _T_2109;	// sequencer-master.scala:273:29, :329:29
      wire _T_2198 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vs2_valid & &tail ?
                io_op_bits_base_vs2_valid : ~(&tail) & _T_2110) : _T_2110;	// sequencer-master.scala:267:35, :273:29, :329:29, util.scala:94:11
      wire _T_2199 = io_op_bits_active_vstx & (_T_291 | _T_132 | _T_4);	// sequencer-master.scala:231:25
      wire _T_2200 = io_op_bits_active_vstx & (_T_292 | _T_133 | _T_5);	// sequencer-master.scala:231:25
      wire _T_2201 = io_op_bits_active_vstx & (_T_293 | _T_134 | _T_6);	// sequencer-master.scala:231:25
      wire _T_2202 = io_op_bits_active_vstx & (_T_294 | _T_135 | _T_7);	// sequencer-master.scala:231:25
      wire _T_2203 = io_op_bits_active_vstx & (_T_295 | _T_136 | _T_8);	// sequencer-master.scala:231:25
      wire _T_2204 = io_op_bits_active_vstx & (_T_296 | _T_137 | _T_9);	// sequencer-master.scala:231:25
      wire _T_2205 = io_op_bits_active_vstx & (_T_297 | _T_138 | _T_10);	// sequencer-master.scala:231:25
      wire _T_2206 = io_op_bits_active_vstx & (&_T_1 | &_T_0 | &tail);	// sequencer-master.scala:231:25, :267:35, util.scala:94:11
      wire _T_2207 = io_op_bits_active_vstx & (_T_291 | _T_132 | _T_4);	// sequencer-master.scala:232:25
      wire _T_2208 = io_op_bits_active_vstx & (_T_292 | _T_133 | _T_5);	// sequencer-master.scala:232:25
      wire _T_2209 = io_op_bits_active_vstx & (_T_293 | _T_134 | _T_6);	// sequencer-master.scala:232:25
      wire _T_2210 = io_op_bits_active_vstx & (_T_294 | _T_135 | _T_7);	// sequencer-master.scala:232:25
      wire _T_2211 = io_op_bits_active_vstx & (_T_295 | _T_136 | _T_8);	// sequencer-master.scala:232:25
      wire _T_2212 = io_op_bits_active_vstx & (_T_296 | _T_137 | _T_9);	// sequencer-master.scala:232:25
      wire _T_2213 = io_op_bits_active_vstx & (_T_297 | _T_138 | _T_10);	// sequencer-master.scala:232:25
      wire _T_2214 = io_op_bits_active_vstx & (&_T_1 | &_T_0 | &tail);	// sequencer-master.scala:232:25, :267:35, util.scala:94:11
      wire _T_2215 = (~io_op_bits_active_vld | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_valid : ~_T_291 & ~_T_132 &
                (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid : ~_T_4 & _T_2191)) :
                _T_2191);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2216 = (~io_op_bits_active_vld | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_valid : ~_T_292 & ~_T_133 &
                (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid : ~_T_5 & _T_2192)) :
                _T_2192);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2217 = (~io_op_bits_active_vld | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_valid : ~_T_293 & ~_T_134 &
                (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid : ~_T_6 & _T_2193)) :
                _T_2193);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2218 = (~io_op_bits_active_vld | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_valid : ~_T_294 & ~_T_135 &
                (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid : ~_T_7 & _T_2194)) :
                _T_2194);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2219 = (~io_op_bits_active_vld | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_valid : ~_T_295 & ~_T_136 &
                (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid : ~_T_8 & _T_2195)) :
                _T_2195);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2220 = (~io_op_bits_active_vld | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_valid : ~_T_296 & ~_T_137 &
                (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid : ~_T_9 & _T_2196)) :
                _T_2196);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2221 = (~io_op_bits_active_vld | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_valid : ~_T_297 & ~_T_138 &
                (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid : ~_T_10 & _T_2197)) :
                _T_2197);	// sequencer-master.scala:273:29, :329:29, :355:25
      wire _T_2222 = (~io_op_bits_active_vld | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vstx ?
                (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_valid : ~(&_T_1) & ~(&_T_0) &
                (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid : ~(&tail) & _T_2198)) :
                _T_2198);	// sequencer-master.scala:267:35, :273:29, :329:29, :355:25, util.scala:94:11
      wire _T_2223 = io_op_bits_active_vld & (_T_291 | _T_132 | _T_4);	// sequencer-master.scala:230:21
      wire _T_2224 = io_op_bits_active_vld & (_T_292 | _T_133 | _T_5);	// sequencer-master.scala:230:21
      wire _T_2225 = io_op_bits_active_vld & (_T_293 | _T_134 | _T_6);	// sequencer-master.scala:230:21
      wire _T_2226 = io_op_bits_active_vld & (_T_294 | _T_135 | _T_7);	// sequencer-master.scala:230:21
      wire _T_2227 = io_op_bits_active_vld & (_T_295 | _T_136 | _T_8);	// sequencer-master.scala:230:21
      wire _T_2228 = io_op_bits_active_vld & (_T_296 | _T_137 | _T_9);	// sequencer-master.scala:230:21
      wire _T_2229 = io_op_bits_active_vld & (_T_297 | _T_138 | _T_10);	// sequencer-master.scala:230:21
      wire _T_2230 = io_op_bits_active_vld & (&_T_1 | &_T_0 | &tail);	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire _T_2231 = _T_3 & (io_op_bits_active_vst | io_op_bits_active_vld | io_op_bits_active_vstx |
                io_op_bits_active_vldx | io_op_bits_active_vamo | io_op_bits_active_vrfirst |
                io_op_bits_active_vrpred | io_op_bits_active_vfconv | io_op_bits_active_vfcmp |
                io_op_bits_active_vfdiv | io_op_bits_active_vfma | io_op_bits_active_vidiv |
                io_op_bits_active_vimul | io_op_bits_active_vipred | io_op_bits_active_vint);	// sequencer-master.scala:265:41
      wire _T_2232 = v_0 & e_0_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2233 = ~e_0_base_vd_pred & e_0_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2234 = ~io_op_bits_base_vp_pred & io_op_bits_base_vp_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2235 = ~e_0_base_vd_pred & ~e_0_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2236 = ~io_op_bits_base_vp_pred & ~io_op_bits_base_vp_scalar;	// types-vxu.scala:119:31, :120:{37,40}
      wire [7:0] _T_2237 = {4'h0, io_op_bits_base_vp_id};	// sequencer-master.scala:141:29, :247:46
      wire _T_2238 = _T_2232 & io_op_bits_base_vp_valid & ~_T_2233 & ~_T_2234 & (_T_2235 & _T_2236 |
                e_0_base_vd_pred & io_op_bits_base_vp_pred) & e_0_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2239 = v_1 & e_1_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2240 = ~e_1_base_vd_pred & e_1_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2241 = ~e_1_base_vd_pred & ~e_1_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2242 = _T_2239 & io_op_bits_base_vp_valid & ~_T_2240 & ~_T_2234 & (_T_2241 & _T_2236 |
                e_1_base_vd_pred & io_op_bits_base_vp_pred) & e_1_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2243 = v_2 & e_2_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2244 = ~e_2_base_vd_pred & e_2_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2245 = ~e_2_base_vd_pred & ~e_2_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2246 = _T_2243 & io_op_bits_base_vp_valid & ~_T_2244 & ~_T_2234 & (_T_2245 & _T_2236 |
                e_2_base_vd_pred & io_op_bits_base_vp_pred) & e_2_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2247 = v_3 & e_3_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2248 = ~e_3_base_vd_pred & e_3_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2249 = ~e_3_base_vd_pred & ~e_3_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2250 = _T_2247 & io_op_bits_base_vp_valid & ~_T_2248 & ~_T_2234 & (_T_2249 & _T_2236 |
                e_3_base_vd_pred & io_op_bits_base_vp_pred) & e_3_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2251 = v_4 & e_4_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2252 = ~e_4_base_vd_pred & e_4_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2253 = ~e_4_base_vd_pred & ~e_4_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2254 = _T_2251 & io_op_bits_base_vp_valid & ~_T_2252 & ~_T_2234 & (_T_2253 & _T_2236 |
                e_4_base_vd_pred & io_op_bits_base_vp_pred) & e_4_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2255 = v_5 & e_5_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2256 = ~e_5_base_vd_pred & e_5_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2257 = ~e_5_base_vd_pred & ~e_5_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2258 = _T_2255 & io_op_bits_base_vp_valid & ~_T_2256 & ~_T_2234 & (_T_2257 & _T_2236 |
                e_5_base_vd_pred & io_op_bits_base_vp_pred) & e_5_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2259 = v_6 & e_6_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2260 = ~e_6_base_vd_pred & e_6_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2261 = ~e_6_base_vd_pred & ~e_6_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2262 = _T_2259 & io_op_bits_base_vp_valid & ~_T_2260 & ~_T_2234 & (_T_2261 & _T_2236 |
                e_6_base_vd_pred & io_op_bits_base_vp_pred) & e_6_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2263 = v_7 & e_7_base_vd_valid;	// sequencer-master.scala:136:44
      wire _T_2264 = ~e_7_base_vd_pred & e_7_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2265 = ~e_7_base_vd_pred & ~e_7_base_vd_scalar;	// types-vxu.scala:119:{31,37}, :120:{37,40}
      wire _T_2266 = _T_2263 & io_op_bits_base_vp_valid & ~_T_2264 & ~_T_2234 & (_T_2265 & _T_2236 |
                e_7_base_vd_pred & io_op_bits_base_vp_pred) & e_7_base_vd_id == _T_2237;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2267 = ~io_op_bits_base_vs1_pred & io_op_bits_base_vs1_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2268 = ~io_op_bits_base_vs1_pred & ~io_op_bits_base_vs1_scalar;	// types-vxu.scala:119:31, :120:{37,40}
      wire _T_2269 = _T_2232 & io_op_bits_base_vs1_valid & ~_T_2233 & ~_T_2267 & (_T_2235 & _T_2268 |
                e_0_base_vd_pred & io_op_bits_base_vs1_pred) & e_0_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2270 = _T_2239 & io_op_bits_base_vs1_valid & ~_T_2240 & ~_T_2267 & (_T_2241 & _T_2268 |
                e_1_base_vd_pred & io_op_bits_base_vs1_pred) & e_1_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2271 = _T_2243 & io_op_bits_base_vs1_valid & ~_T_2244 & ~_T_2267 & (_T_2245 & _T_2268 |
                e_2_base_vd_pred & io_op_bits_base_vs1_pred) & e_2_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2272 = _T_2247 & io_op_bits_base_vs1_valid & ~_T_2248 & ~_T_2267 & (_T_2249 & _T_2268 |
                e_3_base_vd_pred & io_op_bits_base_vs1_pred) & e_3_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2273 = _T_2251 & io_op_bits_base_vs1_valid & ~_T_2252 & ~_T_2267 & (_T_2253 & _T_2268 |
                e_4_base_vd_pred & io_op_bits_base_vs1_pred) & e_4_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2274 = _T_2255 & io_op_bits_base_vs1_valid & ~_T_2256 & ~_T_2267 & (_T_2257 & _T_2268 |
                e_5_base_vd_pred & io_op_bits_base_vs1_pred) & e_5_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2275 = _T_2259 & io_op_bits_base_vs1_valid & ~_T_2260 & ~_T_2267 & (_T_2261 & _T_2268 |
                e_6_base_vd_pred & io_op_bits_base_vs1_pred) & e_6_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2276 = _T_2263 & io_op_bits_base_vs1_valid & ~_T_2264 & ~_T_2267 & (_T_2265 & _T_2268 |
                e_7_base_vd_pred & io_op_bits_base_vs1_pred) & e_7_base_vd_id == io_op_bits_base_vs1_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2277 = ~io_op_bits_base_vs2_pred & io_op_bits_base_vs2_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2278 = ~io_op_bits_base_vs2_pred & ~io_op_bits_base_vs2_scalar;	// types-vxu.scala:119:31, :120:{37,40}
      wire _T_2279 = _T_2232 & io_op_bits_base_vs2_valid & ~_T_2233 & ~_T_2277 & (_T_2235 & _T_2278 |
                e_0_base_vd_pred & io_op_bits_base_vs2_pred) & e_0_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2280 = _T_2239 & io_op_bits_base_vs2_valid & ~_T_2240 & ~_T_2277 & (_T_2241 & _T_2278 |
                e_1_base_vd_pred & io_op_bits_base_vs2_pred) & e_1_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2281 = _T_2243 & io_op_bits_base_vs2_valid & ~_T_2244 & ~_T_2277 & (_T_2245 & _T_2278 |
                e_2_base_vd_pred & io_op_bits_base_vs2_pred) & e_2_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2282 = _T_2247 & io_op_bits_base_vs2_valid & ~_T_2248 & ~_T_2277 & (_T_2249 & _T_2278 |
                e_3_base_vd_pred & io_op_bits_base_vs2_pred) & e_3_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2283 = _T_2251 & io_op_bits_base_vs2_valid & ~_T_2252 & ~_T_2277 & (_T_2253 & _T_2278 |
                e_4_base_vd_pred & io_op_bits_base_vs2_pred) & e_4_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2284 = _T_2255 & io_op_bits_base_vs2_valid & ~_T_2256 & ~_T_2277 & (_T_2257 & _T_2278 |
                e_5_base_vd_pred & io_op_bits_base_vs2_pred) & e_5_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2285 = _T_2259 & io_op_bits_base_vs2_valid & ~_T_2260 & ~_T_2277 & (_T_2261 & _T_2278 |
                e_6_base_vd_pred & io_op_bits_base_vs2_pred) & e_6_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2286 = _T_2263 & io_op_bits_base_vs2_valid & ~_T_2264 & ~_T_2277 & (_T_2265 & _T_2278 |
                e_7_base_vd_pred & io_op_bits_base_vs2_pred) & e_7_base_vd_id == io_op_bits_base_vs2_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2287 = ~io_op_bits_base_vs3_pred & io_op_bits_base_vs3_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2288 = ~io_op_bits_base_vs3_pred & ~io_op_bits_base_vs3_scalar;	// types-vxu.scala:119:31, :120:{37,40}
      wire _T_2289 = _T_2232 & io_op_bits_base_vs3_valid & ~_T_2233 & ~_T_2287 & (_T_2235 & _T_2288 |
                e_0_base_vd_pred & io_op_bits_base_vs3_pred) & e_0_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2290 = _T_2239 & io_op_bits_base_vs3_valid & ~_T_2240 & ~_T_2287 & (_T_2241 & _T_2288 |
                e_1_base_vd_pred & io_op_bits_base_vs3_pred) & e_1_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2291 = _T_2243 & io_op_bits_base_vs3_valid & ~_T_2244 & ~_T_2287 & (_T_2245 & _T_2288 |
                e_2_base_vd_pred & io_op_bits_base_vs3_pred) & e_2_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2292 = _T_2247 & io_op_bits_base_vs3_valid & ~_T_2248 & ~_T_2287 & (_T_2249 & _T_2288 |
                e_3_base_vd_pred & io_op_bits_base_vs3_pred) & e_3_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2293 = _T_2251 & io_op_bits_base_vs3_valid & ~_T_2252 & ~_T_2287 & (_T_2253 & _T_2288 |
                e_4_base_vd_pred & io_op_bits_base_vs3_pred) & e_4_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2294 = _T_2255 & io_op_bits_base_vs3_valid & ~_T_2256 & ~_T_2287 & (_T_2257 & _T_2288 |
                e_5_base_vd_pred & io_op_bits_base_vs3_pred) & e_5_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2295 = _T_2259 & io_op_bits_base_vs3_valid & ~_T_2260 & ~_T_2287 & (_T_2261 & _T_2288 |
                e_6_base_vd_pred & io_op_bits_base_vs3_pred) & e_6_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2296 = _T_2263 & io_op_bits_base_vs3_valid & ~_T_2264 & ~_T_2287 & (_T_2265 & _T_2288 |
                e_7_base_vd_pred & io_op_bits_base_vs3_pred) & e_7_base_vd_id == io_op_bits_base_vs3_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2297 = ~io_op_bits_base_vd_pred & io_op_bits_base_vd_scalar;	// types-vxu.scala:119:{31,37}
      wire _T_2298 = ~io_op_bits_base_vd_pred & ~io_op_bits_base_vd_scalar;	// types-vxu.scala:119:31, :120:{37,40}
      wire _T_2299 = _T_2232 & io_op_bits_base_vd_valid & ~_T_2233 & ~_T_2297 & (_T_2235 & _T_2298 |
                e_0_base_vd_pred & io_op_bits_base_vd_pred) & e_0_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2300 = _T_2239 & io_op_bits_base_vd_valid & ~_T_2240 & ~_T_2297 & (_T_2241 & _T_2298 |
                e_1_base_vd_pred & io_op_bits_base_vd_pred) & e_1_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2301 = _T_2243 & io_op_bits_base_vd_valid & ~_T_2244 & ~_T_2297 & (_T_2245 & _T_2298 |
                e_2_base_vd_pred & io_op_bits_base_vd_pred) & e_2_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2302 = _T_2247 & io_op_bits_base_vd_valid & ~_T_2248 & ~_T_2297 & (_T_2249 & _T_2298 |
                e_3_base_vd_pred & io_op_bits_base_vd_pred) & e_3_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2303 = _T_2251 & io_op_bits_base_vd_valid & ~_T_2252 & ~_T_2297 & (_T_2253 & _T_2298 |
                e_4_base_vd_pred & io_op_bits_base_vd_pred) & e_4_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2304 = _T_2255 & io_op_bits_base_vd_valid & ~_T_2256 & ~_T_2297 & (_T_2257 & _T_2298 |
                e_5_base_vd_pred & io_op_bits_base_vd_pred) & e_5_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2305 = _T_2259 & io_op_bits_base_vd_valid & ~_T_2260 & ~_T_2297 & (_T_2261 & _T_2298 |
                e_6_base_vd_pred & io_op_bits_base_vd_pred) & e_6_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2306 = _T_2263 & io_op_bits_base_vd_valid & ~_T_2264 & ~_T_2297 & (_T_2265 & _T_2298 |
                e_7_base_vd_pred & io_op_bits_base_vd_pred) & e_7_base_vd_id == io_op_bits_base_vd_id;	// sequencer-master.scala:138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, types-vxu.scala:119:31
      wire _T_2307 = ~io_op_bits_base_vd_valid | ~_T_2297 | reset;	// sequencer-master.scala:138:42, :361:{15,16}
      wire _T_2308 = v_0 & e_0_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_0_base_vp_pred &
                e_0_base_vp_scalar) & ~_T_2297 & (~e_0_base_vp_pred & ~e_0_base_vp_scalar & _T_2298 |
                e_0_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_0_base_vp_id} ==
                io_op_bits_base_vd_id | v_0 & e_0_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_0_base_vs1_pred & e_0_base_vs1_scalar) & ~_T_2297 & (~e_0_base_vs1_pred &
                ~e_0_base_vs1_scalar & _T_2298 | e_0_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_0_base_vs1_id == io_op_bits_base_vd_id | v_0 & e_0_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_0_base_vs2_pred & e_0_base_vs2_scalar) & ~_T_2297 &
                (~e_0_base_vs2_pred & ~e_0_base_vs2_scalar & _T_2298 | e_0_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_0_base_vs2_id == io_op_bits_base_vd_id | v_0 &
                e_0_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_0_base_vs3_pred & e_0_base_vs3_scalar)
                & ~_T_2297 & (~e_0_base_vs3_pred & ~e_0_base_vs3_scalar & _T_2298 | e_0_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_0_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2309 = v_1 & e_1_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_1_base_vp_pred &
                e_1_base_vp_scalar) & ~_T_2297 & (~e_1_base_vp_pred & ~e_1_base_vp_scalar & _T_2298 |
                e_1_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_1_base_vp_id} ==
                io_op_bits_base_vd_id | v_1 & e_1_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_1_base_vs1_pred & e_1_base_vs1_scalar) & ~_T_2297 & (~e_1_base_vs1_pred &
                ~e_1_base_vs1_scalar & _T_2298 | e_1_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_1_base_vs1_id == io_op_bits_base_vd_id | v_1 & e_1_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_1_base_vs2_pred & e_1_base_vs2_scalar) & ~_T_2297 &
                (~e_1_base_vs2_pred & ~e_1_base_vs2_scalar & _T_2298 | e_1_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_1_base_vs2_id == io_op_bits_base_vd_id | v_1 &
                e_1_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_1_base_vs3_pred & e_1_base_vs3_scalar)
                & ~_T_2297 & (~e_1_base_vs3_pred & ~e_1_base_vs3_scalar & _T_2298 | e_1_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_1_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2310 = v_2 & e_2_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_2_base_vp_pred &
                e_2_base_vp_scalar) & ~_T_2297 & (~e_2_base_vp_pred & ~e_2_base_vp_scalar & _T_2298 |
                e_2_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_2_base_vp_id} ==
                io_op_bits_base_vd_id | v_2 & e_2_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_2_base_vs1_pred & e_2_base_vs1_scalar) & ~_T_2297 & (~e_2_base_vs1_pred &
                ~e_2_base_vs1_scalar & _T_2298 | e_2_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_2_base_vs1_id == io_op_bits_base_vd_id | v_2 & e_2_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_2_base_vs2_pred & e_2_base_vs2_scalar) & ~_T_2297 &
                (~e_2_base_vs2_pred & ~e_2_base_vs2_scalar & _T_2298 | e_2_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_2_base_vs2_id == io_op_bits_base_vd_id | v_2 &
                e_2_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_2_base_vs3_pred & e_2_base_vs3_scalar)
                & ~_T_2297 & (~e_2_base_vs3_pred & ~e_2_base_vs3_scalar & _T_2298 | e_2_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_2_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2311 = v_3 & e_3_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_3_base_vp_pred &
                e_3_base_vp_scalar) & ~_T_2297 & (~e_3_base_vp_pred & ~e_3_base_vp_scalar & _T_2298 |
                e_3_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_3_base_vp_id} ==
                io_op_bits_base_vd_id | v_3 & e_3_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_3_base_vs1_pred & e_3_base_vs1_scalar) & ~_T_2297 & (~e_3_base_vs1_pred &
                ~e_3_base_vs1_scalar & _T_2298 | e_3_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_3_base_vs1_id == io_op_bits_base_vd_id | v_3 & e_3_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_3_base_vs2_pred & e_3_base_vs2_scalar) & ~_T_2297 &
                (~e_3_base_vs2_pred & ~e_3_base_vs2_scalar & _T_2298 | e_3_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_3_base_vs2_id == io_op_bits_base_vd_id | v_3 &
                e_3_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_3_base_vs3_pred & e_3_base_vs3_scalar)
                & ~_T_2297 & (~e_3_base_vs3_pred & ~e_3_base_vs3_scalar & _T_2298 | e_3_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_3_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2312 = v_4 & e_4_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_4_base_vp_pred &
                e_4_base_vp_scalar) & ~_T_2297 & (~e_4_base_vp_pred & ~e_4_base_vp_scalar & _T_2298 |
                e_4_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_4_base_vp_id} ==
                io_op_bits_base_vd_id | v_4 & e_4_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_4_base_vs1_pred & e_4_base_vs1_scalar) & ~_T_2297 & (~e_4_base_vs1_pred &
                ~e_4_base_vs1_scalar & _T_2298 | e_4_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_4_base_vs1_id == io_op_bits_base_vd_id | v_4 & e_4_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_4_base_vs2_pred & e_4_base_vs2_scalar) & ~_T_2297 &
                (~e_4_base_vs2_pred & ~e_4_base_vs2_scalar & _T_2298 | e_4_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_4_base_vs2_id == io_op_bits_base_vd_id | v_4 &
                e_4_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_4_base_vs3_pred & e_4_base_vs3_scalar)
                & ~_T_2297 & (~e_4_base_vs3_pred & ~e_4_base_vs3_scalar & _T_2298 | e_4_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_4_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2313 = v_5 & e_5_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_5_base_vp_pred &
                e_5_base_vp_scalar) & ~_T_2297 & (~e_5_base_vp_pred & ~e_5_base_vp_scalar & _T_2298 |
                e_5_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_5_base_vp_id} ==
                io_op_bits_base_vd_id | v_5 & e_5_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_5_base_vs1_pred & e_5_base_vs1_scalar) & ~_T_2297 & (~e_5_base_vs1_pred &
                ~e_5_base_vs1_scalar & _T_2298 | e_5_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_5_base_vs1_id == io_op_bits_base_vd_id | v_5 & e_5_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_5_base_vs2_pred & e_5_base_vs2_scalar) & ~_T_2297 &
                (~e_5_base_vs2_pred & ~e_5_base_vs2_scalar & _T_2298 | e_5_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_5_base_vs2_id == io_op_bits_base_vd_id | v_5 &
                e_5_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_5_base_vs3_pred & e_5_base_vs3_scalar)
                & ~_T_2297 & (~e_5_base_vs3_pred & ~e_5_base_vs3_scalar & _T_2298 | e_5_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_5_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2314 = v_6 & e_6_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_6_base_vp_pred &
                e_6_base_vp_scalar) & ~_T_2297 & (~e_6_base_vp_pred & ~e_6_base_vp_scalar & _T_2298 |
                e_6_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_6_base_vp_id} ==
                io_op_bits_base_vd_id | v_6 & e_6_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_6_base_vs1_pred & e_6_base_vs1_scalar) & ~_T_2297 & (~e_6_base_vs1_pred &
                ~e_6_base_vs1_scalar & _T_2298 | e_6_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_6_base_vs1_id == io_op_bits_base_vd_id | v_6 & e_6_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_6_base_vs2_pred & e_6_base_vs2_scalar) & ~_T_2297 &
                (~e_6_base_vs2_pred & ~e_6_base_vs2_scalar & _T_2298 | e_6_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_6_base_vs2_id == io_op_bits_base_vd_id | v_6 &
                e_6_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_6_base_vs3_pred & e_6_base_vs3_scalar)
                & ~_T_2297 & (~e_6_base_vs3_pred & ~e_6_base_vs3_scalar & _T_2298 | e_6_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_6_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2315 = v_7 & e_7_base_vp_valid & io_op_bits_base_vd_valid & ~(~e_7_base_vp_pred &
                e_7_base_vp_scalar) & ~_T_2297 & (~e_7_base_vp_pred & ~e_7_base_vp_scalar & _T_2298 |
                e_7_base_vp_pred & io_op_bits_base_vd_pred) & {4'h0, e_7_base_vp_id} ==
                io_op_bits_base_vd_id | v_7 & e_7_base_vs1_valid & io_op_bits_base_vd_valid &
                ~(~e_7_base_vs1_pred & e_7_base_vs1_scalar) & ~_T_2297 & (~e_7_base_vs1_pred &
                ~e_7_base_vs1_scalar & _T_2298 | e_7_base_vs1_pred & io_op_bits_base_vd_pred) &
                e_7_base_vs1_id == io_op_bits_base_vd_id | v_7 & e_7_base_vs2_valid &
                io_op_bits_base_vd_valid & ~(~e_7_base_vs2_pred & e_7_base_vs2_scalar) & ~_T_2297 &
                (~e_7_base_vs2_pred & ~e_7_base_vs2_scalar & _T_2298 | e_7_base_vs2_pred &
                io_op_bits_base_vd_pred) & e_7_base_vs2_id == io_op_bits_base_vd_id | v_7 &
                e_7_base_vs3_valid & io_op_bits_base_vd_valid & ~(~e_7_base_vs3_pred & e_7_base_vs3_scalar)
                & ~_T_2297 & (~e_7_base_vs3_pred & ~e_7_base_vs3_scalar & _T_2298 | e_7_base_vs3_pred &
                io_op_bits_base_vd_pred) & e_7_base_vs3_id == io_op_bits_base_vd_id;	// sequencer-master.scala:136:44, :138:{11,42}, :139:{39,75}, :140:{37,72}, :141:29, :161:67, :247:46, types-vxu.scala:119:{31,37}, :120:40
      wire _T_2316 = _T_107 | io_op_bits_active_vrpred | io_op_bits_active_vrfirst | reset;	// sequencer-master.scala:298:15
      wire [2:0] _T_2317 = tail - 3'h1;	// util.scala:94:11
      wire _T_2318 = head == 3'h1;	// sequencer-master.scala:267:35, :389:36, :438:21
      wire _T_2319 = head == 3'h2;	// sequencer-master.scala:267:35, :389:36, :438:21
      wire _T_2320 = head == 3'h3;	// sequencer-master.scala:267:35, :389:36, :438:21
      wire _T_2321 = head == 3'h4;	// sequencer-master.scala:389:36, :438:21, util.scala:94:11
      wire _T_2322 = head == 3'h5;	// sequencer-master.scala:183:52, :389:36, :438:21
      wire _T_2323 = head == 3'h6;	// sequencer-master.scala:267:35, :389:36, :438:21
      wire _T_2324 = head == 3'h0;	// sequencer-master.scala:112:17, :372:35, :389:36
      wire _T_2325 = _T_3 & io_op_bits_active_vint & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2326 = _T_3 & io_op_bits_active_vipred & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2327 = _T_3 & io_op_bits_active_vimul & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2328 = _T_400 & ~_T_2316;	// sequencer-master.scala:298:15
      wire _T_2329 = _T_400 & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2330 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2331 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2332 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2333 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2334 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2335 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2336 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2337 = io_op_bits_active_vipred & io_op_bits_base_vs3_valid & _T_2287 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2338 = _T_3 & io_op_bits_active_vfma & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2339 = _T_433 & ~_T_2316;	// sequencer-master.scala:298:15
      wire _T_2340 = _T_433 & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2341 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2342 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2343 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2344 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2345 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2346 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2347 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2348 = io_op_bits_active_vint & io_op_bits_base_vs2_valid & _T_2277 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2349 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_4 | _T_2341 ?
                io_op_bits_sreg_ss2 : e_0_sreg_ss2) : _T_2341 ? io_op_bits_sreg_ss2 : e_0_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2350 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_5 | _T_2342 ?
                io_op_bits_sreg_ss2 : e_1_sreg_ss2) : _T_2342 ? io_op_bits_sreg_ss2 : e_1_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2351 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_6 | _T_2343 ?
                io_op_bits_sreg_ss2 : e_2_sreg_ss2) : _T_2343 ? io_op_bits_sreg_ss2 : e_2_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2352 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_7 | _T_2344 ?
                io_op_bits_sreg_ss2 : e_3_sreg_ss2) : _T_2344 ? io_op_bits_sreg_ss2 : e_3_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2353 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_8 | _T_2345 ?
                io_op_bits_sreg_ss2 : e_4_sreg_ss2) : _T_2345 ? io_op_bits_sreg_ss2 : e_4_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2354 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_9 | _T_2346 ?
                io_op_bits_sreg_ss2 : e_5_sreg_ss2) : _T_2346 ? io_op_bits_sreg_ss2 : e_5_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2355 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (_T_10 | _T_2347 ?
                io_op_bits_sreg_ss2 : e_6_sreg_ss2) : _T_2347 ? io_op_bits_sreg_ss2 : e_6_sreg_ss2;	// sequencer-master.scala:332:31
      wire [63:0] _T_2356 = io_op_bits_active_vipred & io_op_bits_base_vs2_valid & _T_2277 ? (&tail | _T_2348 ?
                io_op_bits_sreg_ss2 : e_7_sreg_ss2) : _T_2348 ? io_op_bits_sreg_ss2 : e_7_sreg_ss2;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2357 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2358 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2359 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2360 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2361 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2362 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2363 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2364 = io_op_bits_active_vimul & io_op_bits_base_vs2_valid & _T_2277 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2365 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_4 | _T_2357 ?
                io_op_bits_sreg_ss2 : _T_2349) : _T_2357 ? io_op_bits_sreg_ss2 : _T_2349;	// sequencer-master.scala:332:31
      wire [63:0] _T_2366 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_5 | _T_2358 ?
                io_op_bits_sreg_ss2 : _T_2350) : _T_2358 ? io_op_bits_sreg_ss2 : _T_2350;	// sequencer-master.scala:332:31
      wire [63:0] _T_2367 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_6 | _T_2359 ?
                io_op_bits_sreg_ss2 : _T_2351) : _T_2359 ? io_op_bits_sreg_ss2 : _T_2351;	// sequencer-master.scala:332:31
      wire [63:0] _T_2368 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_7 | _T_2360 ?
                io_op_bits_sreg_ss2 : _T_2352) : _T_2360 ? io_op_bits_sreg_ss2 : _T_2352;	// sequencer-master.scala:332:31
      wire [63:0] _T_2369 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_8 | _T_2361 ?
                io_op_bits_sreg_ss2 : _T_2353) : _T_2361 ? io_op_bits_sreg_ss2 : _T_2353;	// sequencer-master.scala:332:31
      wire [63:0] _T_2370 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_9 | _T_2362 ?
                io_op_bits_sreg_ss2 : _T_2354) : _T_2362 ? io_op_bits_sreg_ss2 : _T_2354;	// sequencer-master.scala:332:31
      wire [63:0] _T_2371 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_10 | _T_2363 ?
                io_op_bits_sreg_ss2 : _T_2355) : _T_2363 ? io_op_bits_sreg_ss2 : _T_2355;	// sequencer-master.scala:332:31
      wire [63:0] _T_2372 = io_op_bits_active_vidiv & io_op_bits_base_vs2_valid & _T_2277 ? (&tail | _T_2364 ?
                io_op_bits_sreg_ss2 : _T_2356) : _T_2364 ? io_op_bits_sreg_ss2 : _T_2356;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2373 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2374 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2375 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2376 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2377 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2378 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2379 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2380 = io_op_bits_active_vfma & io_op_bits_base_vs2_valid & _T_2277 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2381 = _T_3 & io_op_bits_active_vfcmp & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2382 = _T_3 & io_op_bits_active_vfconv & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2383 = _T_3 & io_op_bits_active_vrpred & ~_T_2316;	// sequencer-master.scala:298:15
      wire _T_2384 = _T_3 & io_op_bits_active_vrfirst & ~_T_2316;	// sequencer-master.scala:298:15
      wire _T_2385 = _T_3 & io_op_bits_active_vamo & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2386 = _T_3 & io_op_bits_active_vldx & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2387 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2388 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2389 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2390 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2391 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2392 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2393 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2394 = io_op_bits_active_vint & io_op_bits_base_vs1_valid & _T_2267 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2395 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_4 | _T_2387 ?
                io_op_bits_sreg_ss1 : e_0_sreg_ss1) : _T_2387 ? io_op_bits_sreg_ss1 : e_0_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2396 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_5 | _T_2388 ?
                io_op_bits_sreg_ss1 : e_1_sreg_ss1) : _T_2388 ? io_op_bits_sreg_ss1 : e_1_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2397 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_6 | _T_2389 ?
                io_op_bits_sreg_ss1 : e_2_sreg_ss1) : _T_2389 ? io_op_bits_sreg_ss1 : e_2_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2398 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_7 | _T_2390 ?
                io_op_bits_sreg_ss1 : e_3_sreg_ss1) : _T_2390 ? io_op_bits_sreg_ss1 : e_3_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2399 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_8 | _T_2391 ?
                io_op_bits_sreg_ss1 : e_4_sreg_ss1) : _T_2391 ? io_op_bits_sreg_ss1 : e_4_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2400 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_9 | _T_2392 ?
                io_op_bits_sreg_ss1 : e_5_sreg_ss1) : _T_2392 ? io_op_bits_sreg_ss1 : e_5_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2401 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (_T_10 | _T_2393 ?
                io_op_bits_sreg_ss1 : e_6_sreg_ss1) : _T_2393 ? io_op_bits_sreg_ss1 : e_6_sreg_ss1;	// sequencer-master.scala:332:31
      wire [63:0] _T_2402 = io_op_bits_active_vipred & io_op_bits_base_vs1_valid & _T_2267 ? (&tail | _T_2394 ?
                io_op_bits_sreg_ss1 : e_7_sreg_ss1) : _T_2394 ? io_op_bits_sreg_ss1 : e_7_sreg_ss1;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2403 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2404 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2405 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2406 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2407 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2408 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2409 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2410 = io_op_bits_active_vimul & io_op_bits_base_vs1_valid & _T_2267 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2411 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_4 | _T_2403 ?
                io_op_bits_sreg_ss1 : _T_2395) : _T_2403 ? io_op_bits_sreg_ss1 : _T_2395;	// sequencer-master.scala:332:31
      wire [63:0] _T_2412 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_5 | _T_2404 ?
                io_op_bits_sreg_ss1 : _T_2396) : _T_2404 ? io_op_bits_sreg_ss1 : _T_2396;	// sequencer-master.scala:332:31
      wire [63:0] _T_2413 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_6 | _T_2405 ?
                io_op_bits_sreg_ss1 : _T_2397) : _T_2405 ? io_op_bits_sreg_ss1 : _T_2397;	// sequencer-master.scala:332:31
      wire [63:0] _T_2414 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_7 | _T_2406 ?
                io_op_bits_sreg_ss1 : _T_2398) : _T_2406 ? io_op_bits_sreg_ss1 : _T_2398;	// sequencer-master.scala:332:31
      wire [63:0] _T_2415 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_8 | _T_2407 ?
                io_op_bits_sreg_ss1 : _T_2399) : _T_2407 ? io_op_bits_sreg_ss1 : _T_2399;	// sequencer-master.scala:332:31
      wire [63:0] _T_2416 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_9 | _T_2408 ?
                io_op_bits_sreg_ss1 : _T_2400) : _T_2408 ? io_op_bits_sreg_ss1 : _T_2400;	// sequencer-master.scala:332:31
      wire [63:0] _T_2417 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_10 | _T_2409 ?
                io_op_bits_sreg_ss1 : _T_2401) : _T_2409 ? io_op_bits_sreg_ss1 : _T_2401;	// sequencer-master.scala:332:31
      wire [63:0] _T_2418 = io_op_bits_active_vidiv & io_op_bits_base_vs1_valid & _T_2267 ? (&tail | _T_2410 ?
                io_op_bits_sreg_ss1 : _T_2402) : _T_2410 ? io_op_bits_sreg_ss1 : _T_2402;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2419 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2420 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2421 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2422 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2423 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2424 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2425 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2426 = io_op_bits_active_vfma & io_op_bits_base_vs1_valid & _T_2267 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2427 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_4 | _T_2419 ?
                io_op_bits_sreg_ss1 : _T_2411) : _T_2419 ? io_op_bits_sreg_ss1 : _T_2411;	// sequencer-master.scala:332:31
      wire [63:0] _T_2428 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_5 | _T_2420 ?
                io_op_bits_sreg_ss1 : _T_2412) : _T_2420 ? io_op_bits_sreg_ss1 : _T_2412;	// sequencer-master.scala:332:31
      wire [63:0] _T_2429 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_6 | _T_2421 ?
                io_op_bits_sreg_ss1 : _T_2413) : _T_2421 ? io_op_bits_sreg_ss1 : _T_2413;	// sequencer-master.scala:332:31
      wire [63:0] _T_2430 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_7 | _T_2422 ?
                io_op_bits_sreg_ss1 : _T_2414) : _T_2422 ? io_op_bits_sreg_ss1 : _T_2414;	// sequencer-master.scala:332:31
      wire [63:0] _T_2431 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_8 | _T_2423 ?
                io_op_bits_sreg_ss1 : _T_2415) : _T_2423 ? io_op_bits_sreg_ss1 : _T_2415;	// sequencer-master.scala:332:31
      wire [63:0] _T_2432 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_9 | _T_2424 ?
                io_op_bits_sreg_ss1 : _T_2416) : _T_2424 ? io_op_bits_sreg_ss1 : _T_2416;	// sequencer-master.scala:332:31
      wire [63:0] _T_2433 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_10 | _T_2425 ?
                io_op_bits_sreg_ss1 : _T_2417) : _T_2425 ? io_op_bits_sreg_ss1 : _T_2417;	// sequencer-master.scala:332:31
      wire [63:0] _T_2434 = io_op_bits_active_vfdiv & io_op_bits_base_vs1_valid & _T_2267 ? (&tail | _T_2426 ?
                io_op_bits_sreg_ss1 : _T_2418) : _T_2426 ? io_op_bits_sreg_ss1 : _T_2418;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2435 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2436 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2437 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2438 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2439 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2440 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2441 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2442 = io_op_bits_active_vfcmp & io_op_bits_base_vs1_valid & _T_2267 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2443 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_4 | _T_2435 ?
                io_op_bits_sreg_ss1 : _T_2427) : _T_2435 ? io_op_bits_sreg_ss1 : _T_2427;	// sequencer-master.scala:332:31
      wire [63:0] _T_2444 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_5 | _T_2436 ?
                io_op_bits_sreg_ss1 : _T_2428) : _T_2436 ? io_op_bits_sreg_ss1 : _T_2428;	// sequencer-master.scala:332:31
      wire [63:0] _T_2445 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_6 | _T_2437 ?
                io_op_bits_sreg_ss1 : _T_2429) : _T_2437 ? io_op_bits_sreg_ss1 : _T_2429;	// sequencer-master.scala:332:31
      wire [63:0] _T_2446 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_7 | _T_2438 ?
                io_op_bits_sreg_ss1 : _T_2430) : _T_2438 ? io_op_bits_sreg_ss1 : _T_2430;	// sequencer-master.scala:332:31
      wire [63:0] _T_2447 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_8 | _T_2439 ?
                io_op_bits_sreg_ss1 : _T_2431) : _T_2439 ? io_op_bits_sreg_ss1 : _T_2431;	// sequencer-master.scala:332:31
      wire [63:0] _T_2448 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_9 | _T_2440 ?
                io_op_bits_sreg_ss1 : _T_2432) : _T_2440 ? io_op_bits_sreg_ss1 : _T_2432;	// sequencer-master.scala:332:31
      wire [63:0] _T_2449 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (_T_10 | _T_2441 ?
                io_op_bits_sreg_ss1 : _T_2433) : _T_2441 ? io_op_bits_sreg_ss1 : _T_2433;	// sequencer-master.scala:332:31
      wire [63:0] _T_2450 = io_op_bits_active_vfconv & io_op_bits_base_vs1_valid & _T_2267 ? (&tail | _T_2442 ?
                io_op_bits_sreg_ss1 : _T_2434) : _T_2442 ? io_op_bits_sreg_ss1 : _T_2434;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2451 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_4;	// sequencer-master.scala:332:31
      wire [63:0] _T_2452 = _T_2451 ? io_op_bits_sreg_ss1 : _T_2443;	// sequencer-master.scala:332:31
      wire _T_2453 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_5;	// sequencer-master.scala:332:31
      wire [63:0] _T_2454 = _T_2453 ? io_op_bits_sreg_ss1 : _T_2444;	// sequencer-master.scala:332:31
      wire _T_2455 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_6;	// sequencer-master.scala:332:31
      wire [63:0] _T_2456 = _T_2455 ? io_op_bits_sreg_ss1 : _T_2445;	// sequencer-master.scala:332:31
      wire _T_2457 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_7;	// sequencer-master.scala:332:31
      wire [63:0] _T_2458 = _T_2457 ? io_op_bits_sreg_ss1 : _T_2446;	// sequencer-master.scala:332:31
      wire _T_2459 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_8;	// sequencer-master.scala:332:31
      wire [63:0] _T_2460 = _T_2459 ? io_op_bits_sreg_ss1 : _T_2447;	// sequencer-master.scala:332:31
      wire _T_2461 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_9;	// sequencer-master.scala:332:31
      wire [63:0] _T_2462 = _T_2461 ? io_op_bits_sreg_ss1 : _T_2448;	// sequencer-master.scala:332:31
      wire _T_2463 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & _T_10;	// sequencer-master.scala:332:31
      wire [63:0] _T_2464 = _T_2463 ? io_op_bits_sreg_ss1 : _T_2449;	// sequencer-master.scala:332:31
      wire _T_2465 = io_op_bits_active_vrfirst & io_op_bits_base_vs1_valid & _T_2267 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire [63:0] _T_2466 = _T_2465 ? io_op_bits_sreg_ss1 : _T_2450;	// sequencer-master.scala:332:31
      wire [63:0] _T_2467 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_291 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_4 | _T_2451 ?
                io_op_bits_sreg_ss1 : _T_2443) : _T_2452) : _T_2452;	// sequencer-master.scala:332:31
      wire [63:0] _T_2468 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_292 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_5 | _T_2453 ?
                io_op_bits_sreg_ss1 : _T_2444) : _T_2454) : _T_2454;	// sequencer-master.scala:332:31
      wire [63:0] _T_2469 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_293 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_6 | _T_2455 ?
                io_op_bits_sreg_ss1 : _T_2445) : _T_2456) : _T_2456;	// sequencer-master.scala:332:31
      wire [63:0] _T_2470 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_294 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_7 | _T_2457 ?
                io_op_bits_sreg_ss1 : _T_2446) : _T_2458) : _T_2458;	// sequencer-master.scala:332:31
      wire [63:0] _T_2471 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_295 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_8 | _T_2459 ?
                io_op_bits_sreg_ss1 : _T_2447) : _T_2460) : _T_2460;	// sequencer-master.scala:332:31
      wire [63:0] _T_2472 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_296 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_9 | _T_2461 ?
                io_op_bits_sreg_ss1 : _T_2448) : _T_2462) : _T_2462;	// sequencer-master.scala:332:31
      wire [63:0] _T_2473 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & _T_297 ?
                io_op_bits_sreg_ss2 : io_op_bits_base_vs1_valid & _T_2267 ? (_T_10 | _T_2463 ?
                io_op_bits_sreg_ss1 : _T_2449) : _T_2464) : _T_2464;	// sequencer-master.scala:332:31
      wire [63:0] _T_2474 = io_op_bits_active_vamo ? (io_op_bits_base_vs2_valid & _T_2277 & &_T_1 ? io_op_bits_sreg_ss2
                : io_op_bits_base_vs1_valid & _T_2267 ? (&tail | _T_2465 ? io_op_bits_sreg_ss1 : _T_2450) :
                _T_2466) : _T_2466;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2475 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_4;	// sequencer-master.scala:332:31
      wire _T_2476 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_5;	// sequencer-master.scala:332:31
      wire _T_2477 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_6;	// sequencer-master.scala:332:31
      wire _T_2478 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_7;	// sequencer-master.scala:332:31
      wire _T_2479 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_8;	// sequencer-master.scala:332:31
      wire _T_2480 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_9;	// sequencer-master.scala:332:31
      wire _T_2481 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & _T_10;	// sequencer-master.scala:332:31
      wire _T_2482 = io_op_bits_active_vldx & io_op_bits_base_vs2_valid & _T_2277 & &tail;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
      wire _T_2483 = _T_3 & io_op_bits_active_vstx & ~_T_2307;	// sequencer-master.scala:353:15, :361:15
      wire _T_2484 = _T_3 & io_op_bits_active_vld & ~_T_2307;	// sequencer-master.scala:361:15
      wire _T_2485 = _T_3 & io_op_bits_active_vst & ~_T_2307;	// sequencer-master.scala:353:15, :361:15
      wire _T_2486 = io_op_bits_base_vs1_valid & _T_2268;	// sequencer-master.scala:218:69
      wire _T_2487 = io_op_bits_base_vs2_valid & _T_2278;	// sequencer-master.scala:218:69
      wire [2:0] _T_2488 = {2'h0, _T_2486} + {1'h0, {1'h0, _T_2487} + {1'h0, io_op_bits_base_vs3_valid & _T_2288}};	// Bitwise.scala:48:55, compatibility.scala:120:12, sequencer-master.scala:218:69, :499:57
      wire [2:0] _T_2489 = |_T_2488 ? _T_2488 : {2'h0, ~io_op_bits_active_vipred};	// sequencer-master.scala:220:21, :222:{12,17}, :499:57
      wire _T_2490 = io_op_bits_base_vd_valid & _T_2298;	// sequencer-master.scala:218:69
      wire [1:0] _T_2491 = _T_2489[1:0];	// sequencer-master.scala:230:21
      wire [3:0] _T_2492 = {1'h0, _T_2489} + 4'h2;	// compatibility.scala:120:12, sequencer-master.scala:247:56, util.scala:94:11
      wire [3:0] _T_2493 = io_op_bits_active_vint ? (_T_2298 ? (_T_4 ? _T_2492 : e_0_wport_sram) : _T_4 ? 4'h0 :
                e_0_wport_sram) : e_0_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2494 = io_op_bits_active_vint ? (_T_2298 ? (_T_5 ? _T_2492 : e_1_wport_sram) : _T_5 ? 4'h0 :
                e_1_wport_sram) : e_1_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2495 = io_op_bits_active_vint ? (_T_2298 ? (_T_6 ? _T_2492 : e_2_wport_sram) : _T_6 ? 4'h0 :
                e_2_wport_sram) : e_2_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2496 = io_op_bits_active_vint ? (_T_2298 ? (_T_7 ? _T_2492 : e_3_wport_sram) : _T_7 ? 4'h0 :
                e_3_wport_sram) : e_3_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2497 = io_op_bits_active_vint ? (_T_2298 ? (_T_8 ? _T_2492 : e_4_wport_sram) : _T_8 ? 4'h0 :
                e_4_wport_sram) : e_4_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2498 = io_op_bits_active_vint ? (_T_2298 ? (_T_9 ? _T_2492 : e_5_wport_sram) : _T_9 ? 4'h0 :
                e_5_wport_sram) : e_5_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2499 = io_op_bits_active_vint ? (_T_2298 ? (_T_10 ? _T_2492 : e_6_wport_sram) : _T_10 ? 4'h0 :
                e_6_wport_sram) : e_6_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2500 = io_op_bits_active_vint ? (_T_2298 ? (&tail ? _T_2492 : e_7_wport_sram) : &tail ? 4'h0 :
                e_7_wport_sram) : e_7_wport_sram;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2501 = _T_2492[2:0];	// sequencer-master.scala:236:63
      wire [2:0] _T_2502 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_4 ? _T_2501 : e_0_wport_pred) :
                _T_4 ? 3'h0 : e_0_wport_pred) : e_0_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2503 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_5 ? _T_2501 : e_1_wport_pred) :
                _T_5 ? 3'h0 : e_1_wport_pred) : e_1_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2504 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_6 ? _T_2501 : e_2_wport_pred) :
                _T_6 ? 3'h0 : e_2_wport_pred) : e_2_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2505 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_7 ? _T_2501 : e_3_wport_pred) :
                _T_7 ? 3'h0 : e_3_wport_pred) : e_3_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2506 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_8 ? _T_2501 : e_4_wport_pred) :
                _T_8 ? 3'h0 : e_4_wport_pred) : e_4_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2507 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_9 ? _T_2501 : e_5_wport_pred) :
                _T_9 ? 3'h0 : e_5_wport_pred) : e_5_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2508 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (_T_10 ? _T_2501 : e_6_wport_pred) :
                _T_10 ? 3'h0 : e_6_wport_pred) : e_6_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2509 = io_op_bits_active_vint ? (io_op_bits_base_vd_pred ? (&tail ? _T_2501 : e_7_wport_pred) :
                &tail ? 3'h0 : e_7_wport_pred) : e_7_wport_pred;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [1:0] _T_2510 = io_op_bits_active_vipred ? (_T_4 | _T_1631 ? _T_2491 : e_0_rports) : _T_1631 ? _T_2491 :
                e_0_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2511 = io_op_bits_active_vipred ? (_T_5 | _T_1632 ? _T_2491 : e_1_rports) : _T_1632 ? _T_2491 :
                e_1_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2512 = io_op_bits_active_vipred ? (_T_6 | _T_1633 ? _T_2491 : e_2_rports) : _T_1633 ? _T_2491 :
                e_2_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2513 = io_op_bits_active_vipred ? (_T_7 | _T_1634 ? _T_2491 : e_3_rports) : _T_1634 ? _T_2491 :
                e_3_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2514 = io_op_bits_active_vipred ? (_T_8 | _T_1635 ? _T_2491 : e_4_rports) : _T_1635 ? _T_2491 :
                e_4_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2515 = io_op_bits_active_vipred ? (_T_9 | _T_1636 ? _T_2491 : e_5_rports) : _T_1636 ? _T_2491 :
                e_5_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2516 = io_op_bits_active_vipred ? (_T_10 | _T_1637 ? _T_2491 : e_6_rports) : _T_1637 ? _T_2491 :
                e_6_rports;	// sequencer-master.scala:230:21
      wire [1:0] _T_2517 = io_op_bits_active_vipred ? (&tail | _T_1638 ? _T_2491 : e_7_rports) : _T_1638 ? _T_2491 :
                e_7_rports;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [3:0] _T_2518 = {1'h0, _T_2489} + 4'h1;	// compatibility.scala:120:12, sequencer-master.scala:247:56, util.scala:94:11
      wire [3:0] _T_2519 = io_op_bits_active_vipred ? (_T_2298 ? (_T_4 ? _T_2518 : _T_2493) : _T_4 ? 4'h0 : _T_2493) :
                _T_2493;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2520 = io_op_bits_active_vipred ? (_T_2298 ? (_T_5 ? _T_2518 : _T_2494) : _T_5 ? 4'h0 : _T_2494) :
                _T_2494;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2521 = io_op_bits_active_vipred ? (_T_2298 ? (_T_6 ? _T_2518 : _T_2495) : _T_6 ? 4'h0 : _T_2495) :
                _T_2495;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2522 = io_op_bits_active_vipred ? (_T_2298 ? (_T_7 ? _T_2518 : _T_2496) : _T_7 ? 4'h0 : _T_2496) :
                _T_2496;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2523 = io_op_bits_active_vipred ? (_T_2298 ? (_T_8 ? _T_2518 : _T_2497) : _T_8 ? 4'h0 : _T_2497) :
                _T_2497;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2524 = io_op_bits_active_vipred ? (_T_2298 ? (_T_9 ? _T_2518 : _T_2498) : _T_9 ? 4'h0 : _T_2498) :
                _T_2498;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2525 = io_op_bits_active_vipred ? (_T_2298 ? (_T_10 ? _T_2518 : _T_2499) : _T_10 ? 4'h0 : _T_2499)
                : _T_2499;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2526 = io_op_bits_active_vipred ? (_T_2298 ? (&tail ? _T_2518 : _T_2500) : &tail ? 4'h0 : _T_2500)
                : _T_2500;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2527 = _T_2518[2:0];	// sequencer-master.scala:236:63
      wire [2:0] _T_2528 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_4 ? _T_2527 : _T_2502) : _T_4 ?
                3'h0 : _T_2502) : _T_2502;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2529 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_5 ? _T_2527 : _T_2503) : _T_5 ?
                3'h0 : _T_2503) : _T_2503;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2530 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_6 ? _T_2527 : _T_2504) : _T_6 ?
                3'h0 : _T_2504) : _T_2504;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2531 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_7 ? _T_2527 : _T_2505) : _T_7 ?
                3'h0 : _T_2505) : _T_2505;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2532 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_8 ? _T_2527 : _T_2506) : _T_8 ?
                3'h0 : _T_2506) : _T_2506;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2533 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_9 ? _T_2527 : _T_2507) : _T_9 ?
                3'h0 : _T_2507) : _T_2507;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2534 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (_T_10 ? _T_2527 : _T_2508) : _T_10 ?
                3'h0 : _T_2508) : _T_2508;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2535 = io_op_bits_active_vipred ? (io_op_bits_base_vd_pred ? (&tail ? _T_2527 : _T_2509) : &tail ?
                3'h0 : _T_2509) : _T_2509;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [3:0] _T_2536 = {1'h0, _T_2489} + 4'h4;	// compatibility.scala:120:12, sequencer-master.scala:247:56, util.scala:94:11
      wire [3:0] _T_2537 = io_op_bits_active_vimul ? (_T_2298 ? (_T_4 ? _T_2536 : _T_2519) : _T_4 ? 4'h0 : _T_2519) :
                _T_2519;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2538 = io_op_bits_active_vimul ? (_T_2298 ? (_T_5 ? _T_2536 : _T_2520) : _T_5 ? 4'h0 : _T_2520) :
                _T_2520;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2539 = io_op_bits_active_vimul ? (_T_2298 ? (_T_6 ? _T_2536 : _T_2521) : _T_6 ? 4'h0 : _T_2521) :
                _T_2521;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2540 = io_op_bits_active_vimul ? (_T_2298 ? (_T_7 ? _T_2536 : _T_2522) : _T_7 ? 4'h0 : _T_2522) :
                _T_2522;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2541 = io_op_bits_active_vimul ? (_T_2298 ? (_T_8 ? _T_2536 : _T_2523) : _T_8 ? 4'h0 : _T_2523) :
                _T_2523;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2542 = io_op_bits_active_vimul ? (_T_2298 ? (_T_9 ? _T_2536 : _T_2524) : _T_9 ? 4'h0 : _T_2524) :
                _T_2524;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2543 = io_op_bits_active_vimul ? (_T_2298 ? (_T_10 ? _T_2536 : _T_2525) : _T_10 ? 4'h0 : _T_2525)
                : _T_2525;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2544 = io_op_bits_active_vimul ? (_T_2298 ? (&tail ? _T_2536 : _T_2526) : &tail ? 4'h0 : _T_2526)
                : _T_2526;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2545 = _T_2536[2:0];	// sequencer-master.scala:236:63
      wire [2:0] _T_2546 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_4 ? _T_2545 : _T_2528) : _T_4 ?
                3'h0 : _T_2528) : _T_2528;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2547 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_5 ? _T_2545 : _T_2529) : _T_5 ?
                3'h0 : _T_2529) : _T_2529;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2548 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_6 ? _T_2545 : _T_2530) : _T_6 ?
                3'h0 : _T_2530) : _T_2530;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2549 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_7 ? _T_2545 : _T_2531) : _T_7 ?
                3'h0 : _T_2531) : _T_2531;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2550 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_8 ? _T_2545 : _T_2532) : _T_8 ?
                3'h0 : _T_2532) : _T_2532;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2551 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_9 ? _T_2545 : _T_2533) : _T_9 ?
                3'h0 : _T_2533) : _T_2533;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2552 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (_T_10 ? _T_2545 : _T_2534) : _T_10 ?
                3'h0 : _T_2534) : _T_2534;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2553 = io_op_bits_active_vimul ? (io_op_bits_base_vd_pred ? (&tail ? _T_2545 : _T_2535) : &tail ?
                3'h0 : _T_2535) : _T_2535;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [1:0] _T_2554 = io_op_bits_active_vidiv ? (_T_132 ? 2'h0 : _T_4 | _T_1719 ? _T_2491 : _T_2510) : _T_1719 ?
                _T_2491 : _T_2510;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2555 = io_op_bits_active_vidiv ? (_T_133 ? 2'h0 : _T_5 | _T_1720 ? _T_2491 : _T_2511) : _T_1720 ?
                _T_2491 : _T_2511;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2556 = io_op_bits_active_vidiv ? (_T_134 ? 2'h0 : _T_6 | _T_1721 ? _T_2491 : _T_2512) : _T_1721 ?
                _T_2491 : _T_2512;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2557 = io_op_bits_active_vidiv ? (_T_135 ? 2'h0 : _T_7 | _T_1722 ? _T_2491 : _T_2513) : _T_1722 ?
                _T_2491 : _T_2513;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2558 = io_op_bits_active_vidiv ? (_T_136 ? 2'h0 : _T_8 | _T_1723 ? _T_2491 : _T_2514) : _T_1723 ?
                _T_2491 : _T_2514;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2559 = io_op_bits_active_vidiv ? (_T_137 ? 2'h0 : _T_9 | _T_1724 ? _T_2491 : _T_2515) : _T_1724 ?
                _T_2491 : _T_2515;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2560 = io_op_bits_active_vidiv ? (_T_138 ? 2'h0 : _T_10 | _T_1725 ? _T_2491 : _T_2516) : _T_1725 ?
                _T_2491 : _T_2516;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2561 = io_op_bits_active_vidiv ? (&_T_0 ? 2'h0 : &tail | _T_1726 ? _T_2491 : _T_2517) : _T_1726 ?
                _T_2491 : _T_2517;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      wire [3:0] _T_2562 = {1'h0, _T_2489} + {1'h0, (_io_op_bits_fn_union_7to6 == 2'h1 ? 3'h5 : 3'h0) |
                {_io_op_bits_fn_union_7to6 == 2'h0 | _io_op_bits_fn_union_7to6 == 2'h2, 2'h0}};	// Mux.scala:19:72, compatibility.scala:120:12, sequencer-master.scala:112:17, :183:52, :247:56, :499:57, types-vxu.scala:53:51, util.scala:94:11
      wire [3:0] _T_2563 = io_op_bits_active_vfma ? (_T_2298 & _T_4 ? _T_2562 : _T_4 | _T_1767 ? 4'h0 : _T_2537) :
                _T_1767 ? 4'h0 : _T_2537;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2564 = io_op_bits_active_vfma ? (_T_2298 & _T_5 ? _T_2562 : _T_5 | _T_1768 ? 4'h0 : _T_2538) :
                _T_1768 ? 4'h0 : _T_2538;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2565 = io_op_bits_active_vfma ? (_T_2298 & _T_6 ? _T_2562 : _T_6 | _T_1769 ? 4'h0 : _T_2539) :
                _T_1769 ? 4'h0 : _T_2539;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2566 = io_op_bits_active_vfma ? (_T_2298 & _T_7 ? _T_2562 : _T_7 | _T_1770 ? 4'h0 : _T_2540) :
                _T_1770 ? 4'h0 : _T_2540;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2567 = io_op_bits_active_vfma ? (_T_2298 & _T_8 ? _T_2562 : _T_8 | _T_1771 ? 4'h0 : _T_2541) :
                _T_1771 ? 4'h0 : _T_2541;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2568 = io_op_bits_active_vfma ? (_T_2298 & _T_9 ? _T_2562 : _T_9 | _T_1772 ? 4'h0 : _T_2542) :
                _T_1772 ? 4'h0 : _T_2542;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2569 = io_op_bits_active_vfma ? (_T_2298 & _T_10 ? _T_2562 : _T_10 | _T_1773 ? 4'h0 : _T_2543) :
                _T_1773 ? 4'h0 : _T_2543;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2570 = io_op_bits_active_vfma ? (_T_2298 & &tail ? _T_2562 : &tail | _T_1774 ? 4'h0 : _T_2544) :
                _T_1774 ? 4'h0 : _T_2544;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2571 = _T_2562[2:0];	// sequencer-master.scala:236:63
      wire [2:0] _T_2572 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_4 ? _T_2571 : _T_4 | _T_1775 ? 3'h0
                : _T_2546) : _T_1775 ? 3'h0 : _T_2546;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2573 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_5 ? _T_2571 : _T_5 | _T_1776 ? 3'h0
                : _T_2547) : _T_1776 ? 3'h0 : _T_2547;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2574 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_6 ? _T_2571 : _T_6 | _T_1777 ? 3'h0
                : _T_2548) : _T_1777 ? 3'h0 : _T_2548;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2575 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_7 ? _T_2571 : _T_7 | _T_1778 ? 3'h0
                : _T_2549) : _T_1778 ? 3'h0 : _T_2549;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2576 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_8 ? _T_2571 : _T_8 | _T_1779 ? 3'h0
                : _T_2550) : _T_1779 ? 3'h0 : _T_2550;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2577 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_9 ? _T_2571 : _T_9 | _T_1780 ? 3'h0
                : _T_2551) : _T_1780 ? 3'h0 : _T_2551;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2578 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & _T_10 ? _T_2571 : _T_10 | _T_1781 ?
                3'h0 : _T_2552) : _T_1781 ? 3'h0 : _T_2552;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2579 = io_op_bits_active_vfma ? (io_op_bits_base_vd_pred & &tail ? _T_2571 : &tail | _T_1782 ?
                3'h0 : _T_2553) : _T_1782 ? 3'h0 : _T_2553;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [1:0] _T_2580 = io_op_bits_active_vfdiv ? (_T_132 ? 2'h0 : _T_4 | _T_1823 ? _T_2491 : _T_2554) : _T_1823 ?
                _T_2491 : _T_2554;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2581 = io_op_bits_active_vfdiv ? (_T_133 ? 2'h0 : _T_5 | _T_1824 ? _T_2491 : _T_2555) : _T_1824 ?
                _T_2491 : _T_2555;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2582 = io_op_bits_active_vfdiv ? (_T_134 ? 2'h0 : _T_6 | _T_1825 ? _T_2491 : _T_2556) : _T_1825 ?
                _T_2491 : _T_2556;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2583 = io_op_bits_active_vfdiv ? (_T_135 ? 2'h0 : _T_7 | _T_1826 ? _T_2491 : _T_2557) : _T_1826 ?
                _T_2491 : _T_2557;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2584 = io_op_bits_active_vfdiv ? (_T_136 ? 2'h0 : _T_8 | _T_1827 ? _T_2491 : _T_2558) : _T_1827 ?
                _T_2491 : _T_2558;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2585 = io_op_bits_active_vfdiv ? (_T_137 ? 2'h0 : _T_9 | _T_1828 ? _T_2491 : _T_2559) : _T_1828 ?
                _T_2491 : _T_2559;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2586 = io_op_bits_active_vfdiv ? (_T_138 ? 2'h0 : _T_10 | _T_1829 ? _T_2491 : _T_2560) : _T_1829 ?
                _T_2491 : _T_2560;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2587 = io_op_bits_active_vfdiv ? (&_T_0 ? 2'h0 : &tail | _T_1830 ? _T_2491 : _T_2561) : _T_1830 ?
                _T_2491 : _T_2561;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      wire [3:0] _T_2588 = io_op_bits_active_vfcmp ? (_T_2298 & _T_4 ? _T_2492 : _T_4 | _T_1871 ? 4'h0 : _T_2563) :
                _T_1871 ? 4'h0 : _T_2563;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2589 = io_op_bits_active_vfcmp ? (_T_2298 & _T_5 ? _T_2492 : _T_5 | _T_1872 ? 4'h0 : _T_2564) :
                _T_1872 ? 4'h0 : _T_2564;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2590 = io_op_bits_active_vfcmp ? (_T_2298 & _T_6 ? _T_2492 : _T_6 | _T_1873 ? 4'h0 : _T_2565) :
                _T_1873 ? 4'h0 : _T_2565;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2591 = io_op_bits_active_vfcmp ? (_T_2298 & _T_7 ? _T_2492 : _T_7 | _T_1874 ? 4'h0 : _T_2566) :
                _T_1874 ? 4'h0 : _T_2566;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2592 = io_op_bits_active_vfcmp ? (_T_2298 & _T_8 ? _T_2492 : _T_8 | _T_1875 ? 4'h0 : _T_2567) :
                _T_1875 ? 4'h0 : _T_2567;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2593 = io_op_bits_active_vfcmp ? (_T_2298 & _T_9 ? _T_2492 : _T_9 | _T_1876 ? 4'h0 : _T_2568) :
                _T_1876 ? 4'h0 : _T_2568;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2594 = io_op_bits_active_vfcmp ? (_T_2298 & _T_10 ? _T_2492 : _T_10 | _T_1877 ? 4'h0 : _T_2569) :
                _T_1877 ? 4'h0 : _T_2569;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2595 = io_op_bits_active_vfcmp ? (_T_2298 & &tail ? _T_2492 : &tail | _T_1878 ? 4'h0 : _T_2570) :
                _T_1878 ? 4'h0 : _T_2570;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2596 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_4 ? _T_2501 : _T_4 | _T_1879 ? 3'h0
                : _T_2572) : _T_1879 ? 3'h0 : _T_2572;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2597 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_5 ? _T_2501 : _T_5 | _T_1880 ? 3'h0
                : _T_2573) : _T_1880 ? 3'h0 : _T_2573;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2598 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_6 ? _T_2501 : _T_6 | _T_1881 ? 3'h0
                : _T_2574) : _T_1881 ? 3'h0 : _T_2574;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2599 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_7 ? _T_2501 : _T_7 | _T_1882 ? 3'h0
                : _T_2575) : _T_1882 ? 3'h0 : _T_2575;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2600 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_8 ? _T_2501 : _T_8 | _T_1883 ? 3'h0
                : _T_2576) : _T_1883 ? 3'h0 : _T_2576;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2601 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_9 ? _T_2501 : _T_9 | _T_1884 ? 3'h0
                : _T_2577) : _T_1884 ? 3'h0 : _T_2577;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2602 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & _T_10 ? _T_2501 : _T_10 | _T_1885 ?
                3'h0 : _T_2578) : _T_1885 ? 3'h0 : _T_2578;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2603 = io_op_bits_active_vfcmp ? (io_op_bits_base_vd_pred & &tail ? _T_2501 : &tail | _T_1886 ?
                3'h0 : _T_2579) : _T_1886 ? 3'h0 : _T_2579;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [1:0] _T_2604 = io_op_bits_active_vfconv ? (_T_4 | _T_1927 ? _T_2491 : _T_2580) : _T_1927 ? _T_2491 :
                _T_2580;	// sequencer-master.scala:230:21
      wire [1:0] _T_2605 = io_op_bits_active_vfconv ? (_T_5 | _T_1928 ? _T_2491 : _T_2581) : _T_1928 ? _T_2491 :
                _T_2581;	// sequencer-master.scala:230:21
      wire [1:0] _T_2606 = io_op_bits_active_vfconv ? (_T_6 | _T_1929 ? _T_2491 : _T_2582) : _T_1929 ? _T_2491 :
                _T_2582;	// sequencer-master.scala:230:21
      wire [1:0] _T_2607 = io_op_bits_active_vfconv ? (_T_7 | _T_1930 ? _T_2491 : _T_2583) : _T_1930 ? _T_2491 :
                _T_2583;	// sequencer-master.scala:230:21
      wire [1:0] _T_2608 = io_op_bits_active_vfconv ? (_T_8 | _T_1931 ? _T_2491 : _T_2584) : _T_1931 ? _T_2491 :
                _T_2584;	// sequencer-master.scala:230:21
      wire [1:0] _T_2609 = io_op_bits_active_vfconv ? (_T_9 | _T_1932 ? _T_2491 : _T_2585) : _T_1932 ? _T_2491 :
                _T_2585;	// sequencer-master.scala:230:21
      wire [1:0] _T_2610 = io_op_bits_active_vfconv ? (_T_10 | _T_1933 ? _T_2491 : _T_2586) : _T_1933 ? _T_2491 :
                _T_2586;	// sequencer-master.scala:230:21
      wire [1:0] _T_2611 = io_op_bits_active_vfconv ? (&tail | _T_1934 ? _T_2491 : _T_2587) : _T_1934 ? _T_2491 :
                _T_2587;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [3:0] _T_2612 = {1'h0, _T_2489} + 4'h3;	// compatibility.scala:120:12, sequencer-master.scala:247:56, util.scala:94:11
      wire [3:0] _T_2613 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_4 ? _T_2612 : _T_2588) : _T_4 ? 4'h0 : _T_2588) :
                _T_2588;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2614 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_5 ? _T_2612 : _T_2589) : _T_5 ? 4'h0 : _T_2589) :
                _T_2589;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2615 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_6 ? _T_2612 : _T_2590) : _T_6 ? 4'h0 : _T_2590) :
                _T_2590;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2616 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_7 ? _T_2612 : _T_2591) : _T_7 ? 4'h0 : _T_2591) :
                _T_2591;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2617 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_8 ? _T_2612 : _T_2592) : _T_8 ? 4'h0 : _T_2592) :
                _T_2592;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2618 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_9 ? _T_2612 : _T_2593) : _T_9 ? 4'h0 : _T_2593) :
                _T_2593;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2619 = io_op_bits_active_vfconv ? (_T_2298 ? (_T_10 ? _T_2612 : _T_2594) : _T_10 ? 4'h0 : _T_2594)
                : _T_2594;	// sequencer-master.scala:231:25, :235:65, :247:46
      wire [3:0] _T_2620 = io_op_bits_active_vfconv ? (_T_2298 ? (&tail ? _T_2612 : _T_2595) : &tail ? 4'h0 : _T_2595)
                : _T_2595;	// sequencer-master.scala:231:25, :235:65, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2621 = _T_2612[2:0];	// sequencer-master.scala:236:63
      wire [2:0] _T_2622 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_4 ? _T_2621 : _T_2596) : _T_4 ?
                3'h0 : _T_2596) : _T_2596;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2623 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_5 ? _T_2621 : _T_2597) : _T_5 ?
                3'h0 : _T_2597) : _T_2597;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2624 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_6 ? _T_2621 : _T_2598) : _T_6 ?
                3'h0 : _T_2598) : _T_2598;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2625 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_7 ? _T_2621 : _T_2599) : _T_7 ?
                3'h0 : _T_2599) : _T_2599;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2626 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_8 ? _T_2621 : _T_2600) : _T_8 ?
                3'h0 : _T_2600) : _T_2600;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2627 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_9 ? _T_2621 : _T_2601) : _T_9 ?
                3'h0 : _T_2601) : _T_2601;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2628 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (_T_10 ? _T_2621 : _T_2602) : _T_10 ?
                3'h0 : _T_2602) : _T_2602;	// sequencer-master.scala:112:17, :232:25, :236:63
      wire [2:0] _T_2629 = io_op_bits_active_vfconv ? (io_op_bits_base_vd_pred ? (&tail ? _T_2621 : _T_2603) : &tail ?
                3'h0 : _T_2603) : _T_2603;	// sequencer-master.scala:112:17, :232:25, :236:63, :267:35, util.scala:94:11
      wire [1:0] _T_2630 = io_op_bits_active_vrfirst ? (_T_4 | _T_1975 ? _T_2491 : _T_2604) : _T_1975 ? _T_2491 :
                _T_2604;	// sequencer-master.scala:230:21
      wire [1:0] _T_2631 = io_op_bits_active_vrfirst ? (_T_5 | _T_1976 ? _T_2491 : _T_2605) : _T_1976 ? _T_2491 :
                _T_2605;	// sequencer-master.scala:230:21
      wire [1:0] _T_2632 = io_op_bits_active_vrfirst ? (_T_6 | _T_1977 ? _T_2491 : _T_2606) : _T_1977 ? _T_2491 :
                _T_2606;	// sequencer-master.scala:230:21
      wire [1:0] _T_2633 = io_op_bits_active_vrfirst ? (_T_7 | _T_1978 ? _T_2491 : _T_2607) : _T_1978 ? _T_2491 :
                _T_2607;	// sequencer-master.scala:230:21
      wire [1:0] _T_2634 = io_op_bits_active_vrfirst ? (_T_8 | _T_1979 ? _T_2491 : _T_2608) : _T_1979 ? _T_2491 :
                _T_2608;	// sequencer-master.scala:230:21
      wire [1:0] _T_2635 = io_op_bits_active_vrfirst ? (_T_9 | _T_1980 ? _T_2491 : _T_2609) : _T_1980 ? _T_2491 :
                _T_2609;	// sequencer-master.scala:230:21
      wire [1:0] _T_2636 = io_op_bits_active_vrfirst ? (_T_10 | _T_1981 ? _T_2491 : _T_2610) : _T_1981 ? _T_2491 :
                _T_2610;	// sequencer-master.scala:230:21
      wire [1:0] _T_2637 = io_op_bits_active_vrfirst ? (&tail | _T_1982 ? _T_2491 : _T_2611) : _T_1982 ? _T_2491 :
                _T_2611;	// sequencer-master.scala:230:21, :267:35, util.scala:94:11
      wire [3:0] _T_2638 = io_op_bits_active_vrfirst ? (_T_4 | _T_1983 ? 4'h0 : _T_2613) : _T_1983 ? 4'h0 : _T_2613;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2639 = io_op_bits_active_vrfirst ? (_T_5 | _T_1984 ? 4'h0 : _T_2614) : _T_1984 ? 4'h0 : _T_2614;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2640 = io_op_bits_active_vrfirst ? (_T_6 | _T_1985 ? 4'h0 : _T_2615) : _T_1985 ? 4'h0 : _T_2615;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2641 = io_op_bits_active_vrfirst ? (_T_7 | _T_1986 ? 4'h0 : _T_2616) : _T_1986 ? 4'h0 : _T_2616;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2642 = io_op_bits_active_vrfirst ? (_T_8 | _T_1987 ? 4'h0 : _T_2617) : _T_1987 ? 4'h0 : _T_2617;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2643 = io_op_bits_active_vrfirst ? (_T_9 | _T_1988 ? 4'h0 : _T_2618) : _T_1988 ? 4'h0 : _T_2618;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2644 = io_op_bits_active_vrfirst ? (_T_10 | _T_1989 ? 4'h0 : _T_2619) : _T_1989 ? 4'h0 : _T_2619;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2645 = io_op_bits_active_vrfirst ? (&tail | _T_1990 ? 4'h0 : _T_2620) : _T_1990 ? 4'h0 : _T_2620;	// sequencer-master.scala:231:25, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2646 = io_op_bits_active_vrfirst ? (_T_4 | _T_1991 ? 3'h0 : _T_2622) : _T_1991 ? 3'h0 : _T_2622;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2647 = io_op_bits_active_vrfirst ? (_T_5 | _T_1992 ? 3'h0 : _T_2623) : _T_1992 ? 3'h0 : _T_2623;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2648 = io_op_bits_active_vrfirst ? (_T_6 | _T_1993 ? 3'h0 : _T_2624) : _T_1993 ? 3'h0 : _T_2624;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2649 = io_op_bits_active_vrfirst ? (_T_7 | _T_1994 ? 3'h0 : _T_2625) : _T_1994 ? 3'h0 : _T_2625;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2650 = io_op_bits_active_vrfirst ? (_T_8 | _T_1995 ? 3'h0 : _T_2626) : _T_1995 ? 3'h0 : _T_2626;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2651 = io_op_bits_active_vrfirst ? (_T_9 | _T_1996 ? 3'h0 : _T_2627) : _T_1996 ? 3'h0 : _T_2627;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2652 = io_op_bits_active_vrfirst ? (_T_10 | _T_1997 ? 3'h0 : _T_2628) : _T_1997 ? 3'h0 : _T_2628;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2653 = io_op_bits_active_vrfirst ? (&tail | _T_1998 ? 3'h0 : _T_2629) : _T_1998 ? 3'h0 : _T_2629;	// sequencer-master.scala:112:17, :232:25, :267:35, util.scala:94:11
      wire [1:0] _T_2654 = {1'h0, _T_2486 ? _T_2486 : ~io_op_bits_active_vipred};	// compatibility.scala:120:12, sequencer-master.scala:220:21, :222:12, :230:21
      wire [1:0] _T_2655 = {1'h0, _T_2487 ? _T_2487 : ~io_op_bits_active_vipred};	// compatibility.scala:120:12, sequencer-master.scala:220:21, :222:12, :230:21
      wire [1:0] _T_2656 = io_op_bits_active_vamo ? (_T_314 ? 2'h0 : _T_291 ? _T_2655 : _T_132 ? 2'h0 : _T_4 ? _T_2654
                : _T_2630) : _T_2630;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2657 = io_op_bits_active_vamo ? (_T_315 ? 2'h0 : _T_292 ? _T_2655 : _T_133 ? 2'h0 : _T_5 ? _T_2654
                : _T_2631) : _T_2631;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2658 = io_op_bits_active_vamo ? (_T_316 ? 2'h0 : _T_293 ? _T_2655 : _T_134 ? 2'h0 : _T_6 ? _T_2654
                : _T_2632) : _T_2632;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2659 = io_op_bits_active_vamo ? (_T_317 ? 2'h0 : _T_294 ? _T_2655 : _T_135 ? 2'h0 : _T_7 ? _T_2654
                : _T_2633) : _T_2633;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2660 = io_op_bits_active_vamo ? (_T_318 ? 2'h0 : _T_295 ? _T_2655 : _T_136 ? 2'h0 : _T_8 ? _T_2654
                : _T_2634) : _T_2634;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2661 = io_op_bits_active_vamo ? (_T_319 ? 2'h0 : _T_296 ? _T_2655 : _T_137 ? 2'h0 : _T_9 ? _T_2654
                : _T_2635) : _T_2635;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2662 = io_op_bits_active_vamo ? (_T_320 ? 2'h0 : _T_297 ? _T_2655 : _T_138 ? 2'h0 : _T_10 ?
                _T_2654 : _T_2636) : _T_2636;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2663 = io_op_bits_active_vamo ? (&_T_2 ? 2'h0 : &_T_1 ? _T_2655 : &_T_0 ? 2'h0 : &tail ? _T_2654 :
                _T_2637) : _T_2637;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      wire [1:0] _T_2664 = io_op_bits_active_vldx ? (_T_291 | _T_132 ? 2'h0 : _T_4 ? _T_2655 : _T_2656) : _T_2656;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2665 = io_op_bits_active_vldx ? (_T_292 | _T_133 ? 2'h0 : _T_5 ? _T_2655 : _T_2657) : _T_2657;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2666 = io_op_bits_active_vldx ? (_T_293 | _T_134 ? 2'h0 : _T_6 ? _T_2655 : _T_2658) : _T_2658;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2667 = io_op_bits_active_vldx ? (_T_294 | _T_135 ? 2'h0 : _T_7 ? _T_2655 : _T_2659) : _T_2659;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2668 = io_op_bits_active_vldx ? (_T_295 | _T_136 ? 2'h0 : _T_8 ? _T_2655 : _T_2660) : _T_2660;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2669 = io_op_bits_active_vldx ? (_T_296 | _T_137 ? 2'h0 : _T_9 ? _T_2655 : _T_2661) : _T_2661;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2670 = io_op_bits_active_vldx ? (_T_297 | _T_138 ? 2'h0 : _T_10 ? _T_2655 : _T_2662) : _T_2662;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2671 = io_op_bits_active_vldx ? (&_T_1 | &_T_0 ? 2'h0 : &tail ? _T_2655 : _T_2663) : _T_2663;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      wire [3:0] _T_2672 = io_op_bits_active_vldx ? (_T_291 | _T_132 | _T_4 | _T_2111 ? 4'h0 : _T_2638) : _T_2111 ?
                4'h0 : _T_2638;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2673 = io_op_bits_active_vldx ? (_T_292 | _T_133 | _T_5 | _T_2112 ? 4'h0 : _T_2639) : _T_2112 ?
                4'h0 : _T_2639;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2674 = io_op_bits_active_vldx ? (_T_293 | _T_134 | _T_6 | _T_2113 ? 4'h0 : _T_2640) : _T_2113 ?
                4'h0 : _T_2640;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2675 = io_op_bits_active_vldx ? (_T_294 | _T_135 | _T_7 | _T_2114 ? 4'h0 : _T_2641) : _T_2114 ?
                4'h0 : _T_2641;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2676 = io_op_bits_active_vldx ? (_T_295 | _T_136 | _T_8 | _T_2115 ? 4'h0 : _T_2642) : _T_2115 ?
                4'h0 : _T_2642;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2677 = io_op_bits_active_vldx ? (_T_296 | _T_137 | _T_9 | _T_2116 ? 4'h0 : _T_2643) : _T_2116 ?
                4'h0 : _T_2643;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2678 = io_op_bits_active_vldx ? (_T_297 | _T_138 | _T_10 | _T_2117 ? 4'h0 : _T_2644) : _T_2117 ?
                4'h0 : _T_2644;	// sequencer-master.scala:231:25, :247:46
      wire [3:0] _T_2679 = io_op_bits_active_vldx ? (&_T_1 | &_T_0 | &tail | _T_2118 ? 4'h0 : _T_2645) : _T_2118 ?
                4'h0 : _T_2645;	// sequencer-master.scala:231:25, :247:46, :267:35, util.scala:94:11
      wire [2:0] _T_2680 = io_op_bits_active_vldx ? (_T_291 | _T_132 | _T_4 | _T_2119 ? 3'h0 : _T_2646) : _T_2119 ?
                3'h0 : _T_2646;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2681 = io_op_bits_active_vldx ? (_T_292 | _T_133 | _T_5 | _T_2120 ? 3'h0 : _T_2647) : _T_2120 ?
                3'h0 : _T_2647;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2682 = io_op_bits_active_vldx ? (_T_293 | _T_134 | _T_6 | _T_2121 ? 3'h0 : _T_2648) : _T_2121 ?
                3'h0 : _T_2648;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2683 = io_op_bits_active_vldx ? (_T_294 | _T_135 | _T_7 | _T_2122 ? 3'h0 : _T_2649) : _T_2122 ?
                3'h0 : _T_2649;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2684 = io_op_bits_active_vldx ? (_T_295 | _T_136 | _T_8 | _T_2123 ? 3'h0 : _T_2650) : _T_2123 ?
                3'h0 : _T_2650;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2685 = io_op_bits_active_vldx ? (_T_296 | _T_137 | _T_9 | _T_2124 ? 3'h0 : _T_2651) : _T_2124 ?
                3'h0 : _T_2651;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2686 = io_op_bits_active_vldx ? (_T_297 | _T_138 | _T_10 | _T_2125 ? 3'h0 : _T_2652) : _T_2125 ?
                3'h0 : _T_2652;	// sequencer-master.scala:112:17, :232:25
      wire [2:0] _T_2687 = io_op_bits_active_vldx ? (&_T_1 | &_T_0 | &tail | _T_2126 ? 3'h0 : _T_2653) : _T_2126 ?
                3'h0 : _T_2653;	// sequencer-master.scala:112:17, :232:25, :267:35, util.scala:94:11
      wire [1:0] _T_2688 = {1'h0, _T_2490 ? _T_2490 : ~io_op_bits_active_vipred};	// compatibility.scala:120:12, sequencer-master.scala:220:21, :222:12, :230:21
      wire [1:0] _T_2689 = io_op_bits_active_vstx ? (_T_291 ? _T_2688 : _T_132 ? 2'h0 : _T_4 ? _T_2655 : _T_2664) :
                _T_2664;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2690 = io_op_bits_active_vstx ? (_T_292 ? _T_2688 : _T_133 ? 2'h0 : _T_5 ? _T_2655 : _T_2665) :
                _T_2665;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2691 = io_op_bits_active_vstx ? (_T_293 ? _T_2688 : _T_134 ? 2'h0 : _T_6 ? _T_2655 : _T_2666) :
                _T_2666;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2692 = io_op_bits_active_vstx ? (_T_294 ? _T_2688 : _T_135 ? 2'h0 : _T_7 ? _T_2655 : _T_2667) :
                _T_2667;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2693 = io_op_bits_active_vstx ? (_T_295 ? _T_2688 : _T_136 ? 2'h0 : _T_8 ? _T_2655 : _T_2668) :
                _T_2668;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2694 = io_op_bits_active_vstx ? (_T_296 ? _T_2688 : _T_137 ? 2'h0 : _T_9 ? _T_2655 : _T_2669) :
                _T_2669;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2695 = io_op_bits_active_vstx ? (_T_297 ? _T_2688 : _T_138 ? 2'h0 : _T_10 ? _T_2655 : _T_2670) :
                _T_2670;	// sequencer-master.scala:230:21, :499:57
      wire [1:0] _T_2696 = io_op_bits_active_vstx ? (&_T_1 ? _T_2688 : &_T_0 ? 2'h0 : &tail ? _T_2655 : _T_2671) :
                _T_2671;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      wire _T_2697 = io_op_bits_active_vint ? _T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 &
                e_0_raw_0 : e_0_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_2698 = io_op_bits_active_vint ? _T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 &
                e_0_raw_1 : e_0_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_2699 = io_op_bits_active_vint ? _T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 &
                e_0_raw_2 : e_0_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_2700 = io_op_bits_active_vint ? _T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 &
                e_0_raw_3 : e_0_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_2701 = io_op_bits_active_vint ? _T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 &
                e_0_raw_4 : e_0_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_2702 = io_op_bits_active_vint ? _T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 &
                e_0_raw_5 : e_0_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_2703 = io_op_bits_active_vint ? _T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 &
                e_0_raw_6 : e_0_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_2704 = io_op_bits_active_vint ? _T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 &
                e_0_raw_7 : e_0_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_2705 = io_op_bits_active_vint ? _T_2308 & _T_4 | ~_T_4 & e_0_war_0 : e_0_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_2706 = io_op_bits_active_vint ? _T_2309 & _T_4 | ~_T_4 & e_0_war_1 : e_0_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_2707 = io_op_bits_active_vint ? _T_2310 & _T_4 | ~_T_4 & e_0_war_2 : e_0_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_2708 = io_op_bits_active_vint ? _T_2311 & _T_4 | ~_T_4 & e_0_war_3 : e_0_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_2709 = io_op_bits_active_vint ? _T_2312 & _T_4 | ~_T_4 & e_0_war_4 : e_0_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_2710 = io_op_bits_active_vint ? _T_2313 & _T_4 | ~_T_4 & e_0_war_5 : e_0_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_2711 = io_op_bits_active_vint ? _T_2314 & _T_4 | ~_T_4 & e_0_war_6 : e_0_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_2712 = io_op_bits_active_vint ? _T_2315 & _T_4 | ~_T_4 & e_0_war_7 : e_0_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_2713 = io_op_bits_active_vint ? _T_2299 & _T_4 | ~_T_4 & e_0_waw_0 : e_0_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_2714 = io_op_bits_active_vint ? _T_2300 & _T_4 | ~_T_4 & e_0_waw_1 : e_0_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_2715 = io_op_bits_active_vint ? _T_2301 & _T_4 | ~_T_4 & e_0_waw_2 : e_0_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_2716 = io_op_bits_active_vint ? _T_2302 & _T_4 | ~_T_4 & e_0_waw_3 : e_0_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_2717 = io_op_bits_active_vint ? _T_2303 & _T_4 | ~_T_4 & e_0_waw_4 : e_0_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_2718 = io_op_bits_active_vint ? _T_2304 & _T_4 | ~_T_4 & e_0_waw_5 : e_0_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_2719 = io_op_bits_active_vint ? _T_2305 & _T_4 | ~_T_4 & e_0_waw_6 : e_0_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_2720 = io_op_bits_active_vint ? _T_2306 & _T_4 | ~_T_4 & e_0_waw_7 : e_0_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_2721 = io_op_bits_active_vipred ? _T_2289 & _T_4 | _T_2279 & _T_4 | _T_2269 & _T_4 | ~_T_4 &
                _T_2697 : _T_2697;	// sequencer-master.scala:131:52, :183:52
      wire _T_2722 = io_op_bits_active_vipred ? _T_2290 & _T_4 | _T_2280 & _T_4 | _T_2270 & _T_4 | ~_T_4 &
                _T_2698 : _T_2698;	// sequencer-master.scala:131:52, :183:52
      wire _T_2723 = io_op_bits_active_vipred ? _T_2291 & _T_4 | _T_2281 & _T_4 | _T_2271 & _T_4 | ~_T_4 &
                _T_2699 : _T_2699;	// sequencer-master.scala:131:52, :183:52
      wire _T_2724 = io_op_bits_active_vipred ? _T_2292 & _T_4 | _T_2282 & _T_4 | _T_2272 & _T_4 | ~_T_4 &
                _T_2700 : _T_2700;	// sequencer-master.scala:131:52, :183:52
      wire _T_2725 = io_op_bits_active_vipred ? _T_2293 & _T_4 | _T_2283 & _T_4 | _T_2273 & _T_4 | ~_T_4 &
                _T_2701 : _T_2701;	// sequencer-master.scala:131:52, :183:52
      wire _T_2726 = io_op_bits_active_vipred ? _T_2294 & _T_4 | _T_2284 & _T_4 | _T_2274 & _T_4 | ~_T_4 &
                _T_2702 : _T_2702;	// sequencer-master.scala:131:52, :183:52
      wire _T_2727 = io_op_bits_active_vipred ? _T_2295 & _T_4 | _T_2285 & _T_4 | _T_2275 & _T_4 | ~_T_4 &
                _T_2703 : _T_2703;	// sequencer-master.scala:131:52, :183:52
      wire _T_2728 = io_op_bits_active_vipred ? _T_2296 & _T_4 | _T_2286 & _T_4 | _T_2276 & _T_4 | ~_T_4 &
                _T_2704 : _T_2704;	// sequencer-master.scala:131:52, :183:52
      wire _T_2729 = io_op_bits_active_vipred ? _T_2308 & _T_4 | ~_T_4 & _T_2705 : _T_2705;	// sequencer-master.scala:132:52, :184:52
      wire _T_2730 = io_op_bits_active_vipred ? _T_2309 & _T_4 | ~_T_4 & _T_2706 : _T_2706;	// sequencer-master.scala:132:52, :184:52
      wire _T_2731 = io_op_bits_active_vipred ? _T_2310 & _T_4 | ~_T_4 & _T_2707 : _T_2707;	// sequencer-master.scala:132:52, :184:52
      wire _T_2732 = io_op_bits_active_vipred ? _T_2311 & _T_4 | ~_T_4 & _T_2708 : _T_2708;	// sequencer-master.scala:132:52, :184:52
      wire _T_2733 = io_op_bits_active_vipred ? _T_2312 & _T_4 | ~_T_4 & _T_2709 : _T_2709;	// sequencer-master.scala:132:52, :184:52
      wire _T_2734 = io_op_bits_active_vipred ? _T_2313 & _T_4 | ~_T_4 & _T_2710 : _T_2710;	// sequencer-master.scala:132:52, :184:52
      wire _T_2735 = io_op_bits_active_vipred ? _T_2314 & _T_4 | ~_T_4 & _T_2711 : _T_2711;	// sequencer-master.scala:132:52, :184:52
      wire _T_2736 = io_op_bits_active_vipred ? _T_2315 & _T_4 | ~_T_4 & _T_2712 : _T_2712;	// sequencer-master.scala:132:52, :184:52
      wire _T_2737 = io_op_bits_active_vipred ? _T_2299 & _T_4 | ~_T_4 & _T_2713 : _T_2713;	// sequencer-master.scala:133:52, :185:52
      wire _T_2738 = io_op_bits_active_vipred ? _T_2300 & _T_4 | ~_T_4 & _T_2714 : _T_2714;	// sequencer-master.scala:133:52, :185:52
      wire _T_2739 = io_op_bits_active_vipred ? _T_2301 & _T_4 | ~_T_4 & _T_2715 : _T_2715;	// sequencer-master.scala:133:52, :185:52
      wire _T_2740 = io_op_bits_active_vipred ? _T_2302 & _T_4 | ~_T_4 & _T_2716 : _T_2716;	// sequencer-master.scala:133:52, :185:52
      wire _T_2741 = io_op_bits_active_vipred ? _T_2303 & _T_4 | ~_T_4 & _T_2717 : _T_2717;	// sequencer-master.scala:133:52, :185:52
      wire _T_2742 = io_op_bits_active_vipred ? _T_2304 & _T_4 | ~_T_4 & _T_2718 : _T_2718;	// sequencer-master.scala:133:52, :185:52
      wire _T_2743 = io_op_bits_active_vipred ? _T_2305 & _T_4 | ~_T_4 & _T_2719 : _T_2719;	// sequencer-master.scala:133:52, :185:52
      wire _T_2744 = io_op_bits_active_vipred ? _T_2306 & _T_4 | ~_T_4 & _T_2720 : _T_2720;	// sequencer-master.scala:133:52, :185:52
      wire _T_2745 = io_op_bits_active_vimul ? _T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 &
                _T_2721 : _T_2721;	// sequencer-master.scala:131:52, :183:52
      wire _T_2746 = io_op_bits_active_vimul ? _T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 &
                _T_2722 : _T_2722;	// sequencer-master.scala:131:52, :183:52
      wire _T_2747 = io_op_bits_active_vimul ? _T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 &
                _T_2723 : _T_2723;	// sequencer-master.scala:131:52, :183:52
      wire _T_2748 = io_op_bits_active_vimul ? _T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 &
                _T_2724 : _T_2724;	// sequencer-master.scala:131:52, :183:52
      wire _T_2749 = io_op_bits_active_vimul ? _T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 &
                _T_2725 : _T_2725;	// sequencer-master.scala:131:52, :183:52
      wire _T_2750 = io_op_bits_active_vimul ? _T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 &
                _T_2726 : _T_2726;	// sequencer-master.scala:131:52, :183:52
      wire _T_2751 = io_op_bits_active_vimul ? _T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 &
                _T_2727 : _T_2727;	// sequencer-master.scala:131:52, :183:52
      wire _T_2752 = io_op_bits_active_vimul ? _T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 &
                _T_2728 : _T_2728;	// sequencer-master.scala:131:52, :183:52
      wire _T_2753 = io_op_bits_active_vimul ? _T_2308 & _T_4 | ~_T_4 & _T_2729 : _T_2729;	// sequencer-master.scala:132:52, :184:52
      wire _T_2754 = io_op_bits_active_vimul ? _T_2309 & _T_4 | ~_T_4 & _T_2730 : _T_2730;	// sequencer-master.scala:132:52, :184:52
      wire _T_2755 = io_op_bits_active_vimul ? _T_2310 & _T_4 | ~_T_4 & _T_2731 : _T_2731;	// sequencer-master.scala:132:52, :184:52
      wire _T_2756 = io_op_bits_active_vimul ? _T_2311 & _T_4 | ~_T_4 & _T_2732 : _T_2732;	// sequencer-master.scala:132:52, :184:52
      wire _T_2757 = io_op_bits_active_vimul ? _T_2312 & _T_4 | ~_T_4 & _T_2733 : _T_2733;	// sequencer-master.scala:132:52, :184:52
      wire _T_2758 = io_op_bits_active_vimul ? _T_2313 & _T_4 | ~_T_4 & _T_2734 : _T_2734;	// sequencer-master.scala:132:52, :184:52
      wire _T_2759 = io_op_bits_active_vimul ? _T_2314 & _T_4 | ~_T_4 & _T_2735 : _T_2735;	// sequencer-master.scala:132:52, :184:52
      wire _T_2760 = io_op_bits_active_vimul ? _T_2315 & _T_4 | ~_T_4 & _T_2736 : _T_2736;	// sequencer-master.scala:132:52, :184:52
      wire _T_2761 = io_op_bits_active_vimul ? _T_2299 & _T_4 | ~_T_4 & _T_2737 : _T_2737;	// sequencer-master.scala:133:52, :185:52
      wire _T_2762 = io_op_bits_active_vimul ? _T_2300 & _T_4 | ~_T_4 & _T_2738 : _T_2738;	// sequencer-master.scala:133:52, :185:52
      wire _T_2763 = io_op_bits_active_vimul ? _T_2301 & _T_4 | ~_T_4 & _T_2739 : _T_2739;	// sequencer-master.scala:133:52, :185:52
      wire _T_2764 = io_op_bits_active_vimul ? _T_2302 & _T_4 | ~_T_4 & _T_2740 : _T_2740;	// sequencer-master.scala:133:52, :185:52
      wire _T_2765 = io_op_bits_active_vimul ? _T_2303 & _T_4 | ~_T_4 & _T_2741 : _T_2741;	// sequencer-master.scala:133:52, :185:52
      wire _T_2766 = io_op_bits_active_vimul ? _T_2304 & _T_4 | ~_T_4 & _T_2742 : _T_2742;	// sequencer-master.scala:133:52, :185:52
      wire _T_2767 = io_op_bits_active_vimul ? _T_2305 & _T_4 | ~_T_4 & _T_2743 : _T_2743;	// sequencer-master.scala:133:52, :185:52
      wire _T_2768 = io_op_bits_active_vimul ? _T_2306 & _T_4 | ~_T_4 & _T_2744 : _T_2744;	// sequencer-master.scala:133:52, :185:52
      wire _T_2769 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4 |
                ~_T_4 & _T_2745) : _T_2745;	// sequencer-master.scala:131:52, :183:52
      wire _T_2770 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4 |
                ~_T_4 & _T_2746) : _T_2746;	// sequencer-master.scala:131:52, :183:52
      wire _T_2771 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4 |
                ~_T_4 & _T_2747) : _T_2747;	// sequencer-master.scala:131:52, :183:52
      wire _T_2772 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4 |
                ~_T_4 & _T_2748) : _T_2748;	// sequencer-master.scala:131:52, :183:52
      wire _T_2773 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4 |
                ~_T_4 & _T_2749) : _T_2749;	// sequencer-master.scala:131:52, :183:52
      wire _T_2774 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4 |
                ~_T_4 & _T_2750) : _T_2750;	// sequencer-master.scala:131:52, :183:52
      wire _T_2775 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4 |
                ~_T_4 & _T_2751) : _T_2751;	// sequencer-master.scala:131:52, :183:52
      wire _T_2776 = io_op_bits_active_vidiv ? ~_T_132 & (_T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4 |
                ~_T_4 & _T_2752) : _T_2752;	// sequencer-master.scala:131:52, :183:52
      wire _T_2777 = io_op_bits_active_vidiv ? _T_2308 & _T_132 | ~_T_132 & (_T_2308 & _T_4 | ~_T_4 & _T_2753) :
                _T_2753;	// sequencer-master.scala:132:52, :184:52
      wire _T_2778 = io_op_bits_active_vidiv ? _T_2309 & _T_132 | ~_T_132 & (_T_2309 & _T_4 | ~_T_4 & _T_2754) :
                _T_2754;	// sequencer-master.scala:132:52, :184:52
      wire _T_2779 = io_op_bits_active_vidiv ? _T_2310 & _T_132 | ~_T_132 & (_T_2310 & _T_4 | ~_T_4 & _T_2755) :
                _T_2755;	// sequencer-master.scala:132:52, :184:52
      wire _T_2780 = io_op_bits_active_vidiv ? _T_2311 & _T_132 | ~_T_132 & (_T_2311 & _T_4 | ~_T_4 & _T_2756) :
                _T_2756;	// sequencer-master.scala:132:52, :184:52
      wire _T_2781 = io_op_bits_active_vidiv ? _T_2312 & _T_132 | ~_T_132 & (_T_2312 & _T_4 | ~_T_4 & _T_2757) :
                _T_2757;	// sequencer-master.scala:132:52, :184:52
      wire _T_2782 = io_op_bits_active_vidiv ? _T_2313 & _T_132 | ~_T_132 & (_T_2313 & _T_4 | ~_T_4 & _T_2758) :
                _T_2758;	// sequencer-master.scala:132:52, :184:52
      wire _T_2783 = io_op_bits_active_vidiv ? _T_2314 & _T_132 | ~_T_132 & (_T_2314 & _T_4 | ~_T_4 & _T_2759) :
                _T_2759;	// sequencer-master.scala:132:52, :184:52
      wire _T_2784 = io_op_bits_active_vidiv ? _T_2315 & _T_132 | ~_T_132 & (_T_2315 & _T_4 | ~_T_4 & _T_2760) :
                _T_2760;	// sequencer-master.scala:132:52, :184:52
      wire _T_2785 = io_op_bits_active_vidiv ? _T_2299 & _T_132 | ~_T_132 & (_T_2299 & _T_4 | ~_T_4 & _T_2761) :
                _T_2761;	// sequencer-master.scala:133:52, :185:52
      wire _T_2786 = io_op_bits_active_vidiv ? _T_2300 & _T_132 | ~_T_132 & (_T_2300 & _T_4 | ~_T_4 & _T_2762) :
                _T_2762;	// sequencer-master.scala:133:52, :185:52
      wire _T_2787 = io_op_bits_active_vidiv ? _T_2301 & _T_132 | ~_T_132 & (_T_2301 & _T_4 | ~_T_4 & _T_2763) :
                _T_2763;	// sequencer-master.scala:133:52, :185:52
      wire _T_2788 = io_op_bits_active_vidiv ? _T_2302 & _T_132 | ~_T_132 & (_T_2302 & _T_4 | ~_T_4 & _T_2764) :
                _T_2764;	// sequencer-master.scala:133:52, :185:52
      wire _T_2789 = io_op_bits_active_vidiv ? _T_2303 & _T_132 | ~_T_132 & (_T_2303 & _T_4 | ~_T_4 & _T_2765) :
                _T_2765;	// sequencer-master.scala:133:52, :185:52
      wire _T_2790 = io_op_bits_active_vidiv ? _T_2304 & _T_132 | ~_T_132 & (_T_2304 & _T_4 | ~_T_4 & _T_2766) :
                _T_2766;	// sequencer-master.scala:133:52, :185:52
      wire _T_2791 = io_op_bits_active_vidiv ? _T_2305 & _T_132 | ~_T_132 & (_T_2305 & _T_4 | ~_T_4 & _T_2767) :
                _T_2767;	// sequencer-master.scala:133:52, :185:52
      wire _T_2792 = io_op_bits_active_vidiv ? _T_2306 & _T_132 | ~_T_132 & (_T_2306 & _T_4 | ~_T_4 & _T_2768) :
                _T_2768;	// sequencer-master.scala:133:52, :185:52
      wire _T_2793 = io_op_bits_active_vfma ? _T_2289 & _T_4 | _T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4
                | ~_T_4 & _T_2769 : _T_2769;	// sequencer-master.scala:131:52, :183:52
      wire _T_2794 = io_op_bits_active_vfma ? _T_2290 & _T_4 | _T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4
                | ~_T_4 & _T_2770 : _T_2770;	// sequencer-master.scala:131:52, :183:52
      wire _T_2795 = io_op_bits_active_vfma ? _T_2291 & _T_4 | _T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4
                | ~_T_4 & _T_2771 : _T_2771;	// sequencer-master.scala:131:52, :183:52
      wire _T_2796 = io_op_bits_active_vfma ? _T_2292 & _T_4 | _T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4
                | ~_T_4 & _T_2772 : _T_2772;	// sequencer-master.scala:131:52, :183:52
      wire _T_2797 = io_op_bits_active_vfma ? _T_2293 & _T_4 | _T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4
                | ~_T_4 & _T_2773 : _T_2773;	// sequencer-master.scala:131:52, :183:52
      wire _T_2798 = io_op_bits_active_vfma ? _T_2294 & _T_4 | _T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4
                | ~_T_4 & _T_2774 : _T_2774;	// sequencer-master.scala:131:52, :183:52
      wire _T_2799 = io_op_bits_active_vfma ? _T_2295 & _T_4 | _T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4
                | ~_T_4 & _T_2775 : _T_2775;	// sequencer-master.scala:131:52, :183:52
      wire _T_2800 = io_op_bits_active_vfma ? _T_2296 & _T_4 | _T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4
                | ~_T_4 & _T_2776 : _T_2776;	// sequencer-master.scala:131:52, :183:52
      wire _T_2801 = io_op_bits_active_vfma ? _T_2308 & _T_4 | ~_T_4 & _T_2777 : _T_2777;	// sequencer-master.scala:132:52, :184:52
      wire _T_2802 = io_op_bits_active_vfma ? _T_2309 & _T_4 | ~_T_4 & _T_2778 : _T_2778;	// sequencer-master.scala:132:52, :184:52
      wire _T_2803 = io_op_bits_active_vfma ? _T_2310 & _T_4 | ~_T_4 & _T_2779 : _T_2779;	// sequencer-master.scala:132:52, :184:52
      wire _T_2804 = io_op_bits_active_vfma ? _T_2311 & _T_4 | ~_T_4 & _T_2780 : _T_2780;	// sequencer-master.scala:132:52, :184:52
      wire _T_2805 = io_op_bits_active_vfma ? _T_2312 & _T_4 | ~_T_4 & _T_2781 : _T_2781;	// sequencer-master.scala:132:52, :184:52
      wire _T_2806 = io_op_bits_active_vfma ? _T_2313 & _T_4 | ~_T_4 & _T_2782 : _T_2782;	// sequencer-master.scala:132:52, :184:52
      wire _T_2807 = io_op_bits_active_vfma ? _T_2314 & _T_4 | ~_T_4 & _T_2783 : _T_2783;	// sequencer-master.scala:132:52, :184:52
      wire _T_2808 = io_op_bits_active_vfma ? _T_2315 & _T_4 | ~_T_4 & _T_2784 : _T_2784;	// sequencer-master.scala:132:52, :184:52
      wire _T_2809 = io_op_bits_active_vfma ? _T_2299 & _T_4 | ~_T_4 & _T_2785 : _T_2785;	// sequencer-master.scala:133:52, :185:52
      wire _T_2810 = io_op_bits_active_vfma ? _T_2300 & _T_4 | ~_T_4 & _T_2786 : _T_2786;	// sequencer-master.scala:133:52, :185:52
      wire _T_2811 = io_op_bits_active_vfma ? _T_2301 & _T_4 | ~_T_4 & _T_2787 : _T_2787;	// sequencer-master.scala:133:52, :185:52
      wire _T_2812 = io_op_bits_active_vfma ? _T_2302 & _T_4 | ~_T_4 & _T_2788 : _T_2788;	// sequencer-master.scala:133:52, :185:52
      wire _T_2813 = io_op_bits_active_vfma ? _T_2303 & _T_4 | ~_T_4 & _T_2789 : _T_2789;	// sequencer-master.scala:133:52, :185:52
      wire _T_2814 = io_op_bits_active_vfma ? _T_2304 & _T_4 | ~_T_4 & _T_2790 : _T_2790;	// sequencer-master.scala:133:52, :185:52
      wire _T_2815 = io_op_bits_active_vfma ? _T_2305 & _T_4 | ~_T_4 & _T_2791 : _T_2791;	// sequencer-master.scala:133:52, :185:52
      wire _T_2816 = io_op_bits_active_vfma ? _T_2306 & _T_4 | ~_T_4 & _T_2792 : _T_2792;	// sequencer-master.scala:133:52, :185:52
      wire _T_2817 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4 |
                ~_T_4 & _T_2793) : _T_2793;	// sequencer-master.scala:131:52, :183:52
      wire _T_2818 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4 |
                ~_T_4 & _T_2794) : _T_2794;	// sequencer-master.scala:131:52, :183:52
      wire _T_2819 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4 |
                ~_T_4 & _T_2795) : _T_2795;	// sequencer-master.scala:131:52, :183:52
      wire _T_2820 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4 |
                ~_T_4 & _T_2796) : _T_2796;	// sequencer-master.scala:131:52, :183:52
      wire _T_2821 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4 |
                ~_T_4 & _T_2797) : _T_2797;	// sequencer-master.scala:131:52, :183:52
      wire _T_2822 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4 |
                ~_T_4 & _T_2798) : _T_2798;	// sequencer-master.scala:131:52, :183:52
      wire _T_2823 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4 |
                ~_T_4 & _T_2799) : _T_2799;	// sequencer-master.scala:131:52, :183:52
      wire _T_2824 = io_op_bits_active_vfdiv ? ~_T_132 & (_T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4 |
                ~_T_4 & _T_2800) : _T_2800;	// sequencer-master.scala:131:52, :183:52
      wire _T_2825 = io_op_bits_active_vfdiv ? _T_2308 & _T_132 | ~_T_132 & (_T_2308 & _T_4 | ~_T_4 & _T_2801) :
                _T_2801;	// sequencer-master.scala:132:52, :184:52
      wire _T_2826 = io_op_bits_active_vfdiv ? _T_2309 & _T_132 | ~_T_132 & (_T_2309 & _T_4 | ~_T_4 & _T_2802) :
                _T_2802;	// sequencer-master.scala:132:52, :184:52
      wire _T_2827 = io_op_bits_active_vfdiv ? _T_2310 & _T_132 | ~_T_132 & (_T_2310 & _T_4 | ~_T_4 & _T_2803) :
                _T_2803;	// sequencer-master.scala:132:52, :184:52
      wire _T_2828 = io_op_bits_active_vfdiv ? _T_2311 & _T_132 | ~_T_132 & (_T_2311 & _T_4 | ~_T_4 & _T_2804) :
                _T_2804;	// sequencer-master.scala:132:52, :184:52
      wire _T_2829 = io_op_bits_active_vfdiv ? _T_2312 & _T_132 | ~_T_132 & (_T_2312 & _T_4 | ~_T_4 & _T_2805) :
                _T_2805;	// sequencer-master.scala:132:52, :184:52
      wire _T_2830 = io_op_bits_active_vfdiv ? _T_2313 & _T_132 | ~_T_132 & (_T_2313 & _T_4 | ~_T_4 & _T_2806) :
                _T_2806;	// sequencer-master.scala:132:52, :184:52
      wire _T_2831 = io_op_bits_active_vfdiv ? _T_2314 & _T_132 | ~_T_132 & (_T_2314 & _T_4 | ~_T_4 & _T_2807) :
                _T_2807;	// sequencer-master.scala:132:52, :184:52
      wire _T_2832 = io_op_bits_active_vfdiv ? _T_2315 & _T_132 | ~_T_132 & (_T_2315 & _T_4 | ~_T_4 & _T_2808) :
                _T_2808;	// sequencer-master.scala:132:52, :184:52
      wire _T_2833 = io_op_bits_active_vfdiv ? _T_2299 & _T_132 | ~_T_132 & (_T_2299 & _T_4 | ~_T_4 & _T_2809) :
                _T_2809;	// sequencer-master.scala:133:52, :185:52
      wire _T_2834 = io_op_bits_active_vfdiv ? _T_2300 & _T_132 | ~_T_132 & (_T_2300 & _T_4 | ~_T_4 & _T_2810) :
                _T_2810;	// sequencer-master.scala:133:52, :185:52
      wire _T_2835 = io_op_bits_active_vfdiv ? _T_2301 & _T_132 | ~_T_132 & (_T_2301 & _T_4 | ~_T_4 & _T_2811) :
                _T_2811;	// sequencer-master.scala:133:52, :185:52
      wire _T_2836 = io_op_bits_active_vfdiv ? _T_2302 & _T_132 | ~_T_132 & (_T_2302 & _T_4 | ~_T_4 & _T_2812) :
                _T_2812;	// sequencer-master.scala:133:52, :185:52
      wire _T_2837 = io_op_bits_active_vfdiv ? _T_2303 & _T_132 | ~_T_132 & (_T_2303 & _T_4 | ~_T_4 & _T_2813) :
                _T_2813;	// sequencer-master.scala:133:52, :185:52
      wire _T_2838 = io_op_bits_active_vfdiv ? _T_2304 & _T_132 | ~_T_132 & (_T_2304 & _T_4 | ~_T_4 & _T_2814) :
                _T_2814;	// sequencer-master.scala:133:52, :185:52
      wire _T_2839 = io_op_bits_active_vfdiv ? _T_2305 & _T_132 | ~_T_132 & (_T_2305 & _T_4 | ~_T_4 & _T_2815) :
                _T_2815;	// sequencer-master.scala:133:52, :185:52
      wire _T_2840 = io_op_bits_active_vfdiv ? _T_2306 & _T_132 | ~_T_132 & (_T_2306 & _T_4 | ~_T_4 & _T_2816) :
                _T_2816;	// sequencer-master.scala:133:52, :185:52
      wire _T_2841 = io_op_bits_active_vfcmp ? _T_2279 & _T_4 | _T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 &
                _T_2817 : _T_2817;	// sequencer-master.scala:131:52, :183:52
      wire _T_2842 = io_op_bits_active_vfcmp ? _T_2280 & _T_4 | _T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 &
                _T_2818 : _T_2818;	// sequencer-master.scala:131:52, :183:52
      wire _T_2843 = io_op_bits_active_vfcmp ? _T_2281 & _T_4 | _T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 &
                _T_2819 : _T_2819;	// sequencer-master.scala:131:52, :183:52
      wire _T_2844 = io_op_bits_active_vfcmp ? _T_2282 & _T_4 | _T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 &
                _T_2820 : _T_2820;	// sequencer-master.scala:131:52, :183:52
      wire _T_2845 = io_op_bits_active_vfcmp ? _T_2283 & _T_4 | _T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 &
                _T_2821 : _T_2821;	// sequencer-master.scala:131:52, :183:52
      wire _T_2846 = io_op_bits_active_vfcmp ? _T_2284 & _T_4 | _T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 &
                _T_2822 : _T_2822;	// sequencer-master.scala:131:52, :183:52
      wire _T_2847 = io_op_bits_active_vfcmp ? _T_2285 & _T_4 | _T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 &
                _T_2823 : _T_2823;	// sequencer-master.scala:131:52, :183:52
      wire _T_2848 = io_op_bits_active_vfcmp ? _T_2286 & _T_4 | _T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 &
                _T_2824 : _T_2824;	// sequencer-master.scala:131:52, :183:52
      wire _T_2849 = io_op_bits_active_vfcmp ? _T_2308 & _T_4 | ~_T_4 & _T_2825 : _T_2825;	// sequencer-master.scala:132:52, :184:52
      wire _T_2850 = io_op_bits_active_vfcmp ? _T_2309 & _T_4 | ~_T_4 & _T_2826 : _T_2826;	// sequencer-master.scala:132:52, :184:52
      wire _T_2851 = io_op_bits_active_vfcmp ? _T_2310 & _T_4 | ~_T_4 & _T_2827 : _T_2827;	// sequencer-master.scala:132:52, :184:52
      wire _T_2852 = io_op_bits_active_vfcmp ? _T_2311 & _T_4 | ~_T_4 & _T_2828 : _T_2828;	// sequencer-master.scala:132:52, :184:52
      wire _T_2853 = io_op_bits_active_vfcmp ? _T_2312 & _T_4 | ~_T_4 & _T_2829 : _T_2829;	// sequencer-master.scala:132:52, :184:52
      wire _T_2854 = io_op_bits_active_vfcmp ? _T_2313 & _T_4 | ~_T_4 & _T_2830 : _T_2830;	// sequencer-master.scala:132:52, :184:52
      wire _T_2855 = io_op_bits_active_vfcmp ? _T_2314 & _T_4 | ~_T_4 & _T_2831 : _T_2831;	// sequencer-master.scala:132:52, :184:52
      wire _T_2856 = io_op_bits_active_vfcmp ? _T_2315 & _T_4 | ~_T_4 & _T_2832 : _T_2832;	// sequencer-master.scala:132:52, :184:52
      wire _T_2857 = io_op_bits_active_vfcmp ? _T_2299 & _T_4 | ~_T_4 & _T_2833 : _T_2833;	// sequencer-master.scala:133:52, :185:52
      wire _T_2858 = io_op_bits_active_vfcmp ? _T_2300 & _T_4 | ~_T_4 & _T_2834 : _T_2834;	// sequencer-master.scala:133:52, :185:52
      wire _T_2859 = io_op_bits_active_vfcmp ? _T_2301 & _T_4 | ~_T_4 & _T_2835 : _T_2835;	// sequencer-master.scala:133:52, :185:52
      wire _T_2860 = io_op_bits_active_vfcmp ? _T_2302 & _T_4 | ~_T_4 & _T_2836 : _T_2836;	// sequencer-master.scala:133:52, :185:52
      wire _T_2861 = io_op_bits_active_vfcmp ? _T_2303 & _T_4 | ~_T_4 & _T_2837 : _T_2837;	// sequencer-master.scala:133:52, :185:52
      wire _T_2862 = io_op_bits_active_vfcmp ? _T_2304 & _T_4 | ~_T_4 & _T_2838 : _T_2838;	// sequencer-master.scala:133:52, :185:52
      wire _T_2863 = io_op_bits_active_vfcmp ? _T_2305 & _T_4 | ~_T_4 & _T_2839 : _T_2839;	// sequencer-master.scala:133:52, :185:52
      wire _T_2864 = io_op_bits_active_vfcmp ? _T_2306 & _T_4 | ~_T_4 & _T_2840 : _T_2840;	// sequencer-master.scala:133:52, :185:52
      wire _T_2865 = io_op_bits_active_vfconv ? _T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 & _T_2841 : _T_2841;	// sequencer-master.scala:131:52, :183:52
      wire _T_2866 = io_op_bits_active_vfconv ? _T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 & _T_2842 : _T_2842;	// sequencer-master.scala:131:52, :183:52
      wire _T_2867 = io_op_bits_active_vfconv ? _T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 & _T_2843 : _T_2843;	// sequencer-master.scala:131:52, :183:52
      wire _T_2868 = io_op_bits_active_vfconv ? _T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 & _T_2844 : _T_2844;	// sequencer-master.scala:131:52, :183:52
      wire _T_2869 = io_op_bits_active_vfconv ? _T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 & _T_2845 : _T_2845;	// sequencer-master.scala:131:52, :183:52
      wire _T_2870 = io_op_bits_active_vfconv ? _T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 & _T_2846 : _T_2846;	// sequencer-master.scala:131:52, :183:52
      wire _T_2871 = io_op_bits_active_vfconv ? _T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 & _T_2847 : _T_2847;	// sequencer-master.scala:131:52, :183:52
      wire _T_2872 = io_op_bits_active_vfconv ? _T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 & _T_2848 : _T_2848;	// sequencer-master.scala:131:52, :183:52
      wire _T_2873 = io_op_bits_active_vrpred ? _T_2238 & _T_4 | ~_T_4 & _T_2865 : _T_2865;	// sequencer-master.scala:131:52, :183:52
      wire _T_2874 = io_op_bits_active_vrpred ? _T_2242 & _T_4 | ~_T_4 & _T_2866 : _T_2866;	// sequencer-master.scala:131:52, :183:52
      wire _T_2875 = io_op_bits_active_vrpred ? _T_2246 & _T_4 | ~_T_4 & _T_2867 : _T_2867;	// sequencer-master.scala:131:52, :183:52
      wire _T_2876 = io_op_bits_active_vrpred ? _T_2250 & _T_4 | ~_T_4 & _T_2868 : _T_2868;	// sequencer-master.scala:131:52, :183:52
      wire _T_2877 = io_op_bits_active_vrpred ? _T_2254 & _T_4 | ~_T_4 & _T_2869 : _T_2869;	// sequencer-master.scala:131:52, :183:52
      wire _T_2878 = io_op_bits_active_vrpred ? _T_2258 & _T_4 | ~_T_4 & _T_2870 : _T_2870;	// sequencer-master.scala:131:52, :183:52
      wire _T_2879 = io_op_bits_active_vrpred ? _T_2262 & _T_4 | ~_T_4 & _T_2871 : _T_2871;	// sequencer-master.scala:131:52, :183:52
      wire _T_2880 = io_op_bits_active_vrpred ? _T_2266 & _T_4 | ~_T_4 & _T_2872 : _T_2872;	// sequencer-master.scala:131:52, :183:52
      wire _T_2881 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_4 | ~_T_4 & _T_2849 : _T_2849);	// sequencer-master.scala:132:52, :184:52
      wire _T_2882 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_4 | ~_T_4 & _T_2857 : _T_2857);	// sequencer-master.scala:133:52, :185:52
      wire _T_2883 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_4 | ~_T_4 & _T_2850 : _T_2850);	// sequencer-master.scala:132:52, :184:52
      wire _T_2884 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_4 | ~_T_4 & _T_2858 : _T_2858);	// sequencer-master.scala:133:52, :185:52
      wire _T_2885 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_4 | ~_T_4 & _T_2851 : _T_2851);	// sequencer-master.scala:132:52, :184:52
      wire _T_2886 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_4 | ~_T_4 & _T_2859 : _T_2859);	// sequencer-master.scala:133:52, :185:52
      wire _T_2887 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_4 | ~_T_4 & _T_2852 : _T_2852);	// sequencer-master.scala:132:52, :184:52
      wire _T_2888 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_4 | ~_T_4 & _T_2860 : _T_2860);	// sequencer-master.scala:133:52, :185:52
      wire _T_2889 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_4 | ~_T_4 & _T_2853 : _T_2853);	// sequencer-master.scala:132:52, :184:52
      wire _T_2890 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_4 | ~_T_4 & _T_2861 : _T_2861);	// sequencer-master.scala:133:52, :185:52
      wire _T_2891 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_4 | ~_T_4 & _T_2854 : _T_2854);	// sequencer-master.scala:132:52, :184:52
      wire _T_2892 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_4 | ~_T_4 & _T_2862 : _T_2862);	// sequencer-master.scala:133:52, :185:52
      wire _T_2893 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_4 | ~_T_4 & _T_2855 : _T_2855);	// sequencer-master.scala:132:52, :184:52
      wire _T_2894 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_4 | ~_T_4 & _T_2863 : _T_2863);	// sequencer-master.scala:133:52, :185:52
      wire _T_2895 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_4 | ~_T_4 & _T_2856 : _T_2856);	// sequencer-master.scala:132:52, :184:52
      wire _T_2896 = (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_4 | ~_T_4 & _T_2864 : _T_2864);	// sequencer-master.scala:133:52, :185:52
      wire _T_2897 = io_op_bits_active_vrfirst ? _T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 & _T_2873 : _T_2873;	// sequencer-master.scala:131:52, :183:52
      wire _T_2898 = io_op_bits_active_vrfirst ? _T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 & _T_2874 : _T_2874;	// sequencer-master.scala:131:52, :183:52
      wire _T_2899 = io_op_bits_active_vrfirst ? _T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 & _T_2875 : _T_2875;	// sequencer-master.scala:131:52, :183:52
      wire _T_2900 = io_op_bits_active_vrfirst ? _T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 & _T_2876 : _T_2876;	// sequencer-master.scala:131:52, :183:52
      wire _T_2901 = io_op_bits_active_vrfirst ? _T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 & _T_2877 : _T_2877;	// sequencer-master.scala:131:52, :183:52
      wire _T_2902 = io_op_bits_active_vrfirst ? _T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 & _T_2878 : _T_2878;	// sequencer-master.scala:131:52, :183:52
      wire _T_2903 = io_op_bits_active_vrfirst ? _T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 & _T_2879 : _T_2879;	// sequencer-master.scala:131:52, :183:52
      wire _T_2904 = io_op_bits_active_vrfirst ? _T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 & _T_2880 : _T_2880;	// sequencer-master.scala:131:52, :183:52
      wire _T_2905 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_132 | _T_2279 & _T_291 | _T_2238 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2269 & _T_4 | _T_2238 & _T_4 | ~_T_4 & _T_2897)) : _T_2897;	// sequencer-master.scala:131:52, :183:52
      wire _T_2906 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_133 | _T_2280 & _T_291 | _T_2242 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2270 & _T_4 | _T_2242 & _T_4 | ~_T_4 & _T_2898)) : _T_2898;	// sequencer-master.scala:131:52, :183:52
      wire _T_2907 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_134 | _T_2281 & _T_291 | _T_2246 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2271 & _T_4 | _T_2246 & _T_4 | ~_T_4 & _T_2899)) : _T_2899;	// sequencer-master.scala:131:52, :183:52
      wire _T_2908 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_135 | _T_2282 & _T_291 | _T_2250 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2272 & _T_4 | _T_2250 & _T_4 | ~_T_4 & _T_2900)) : _T_2900;	// sequencer-master.scala:131:52, :183:52
      wire _T_2909 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_136 | _T_2283 & _T_291 | _T_2254 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2273 & _T_4 | _T_2254 & _T_4 | ~_T_4 & _T_2901)) : _T_2901;	// sequencer-master.scala:131:52, :183:52
      wire _T_2910 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_137 | _T_2284 & _T_291 | _T_2258 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2274 & _T_4 | _T_2258 & _T_4 | ~_T_4 & _T_2902)) : _T_2902;	// sequencer-master.scala:131:52, :183:52
      wire _T_2911 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & _T_138 | _T_2285 & _T_291 | _T_2262 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2275 & _T_4 | _T_2262 & _T_4 | ~_T_4 & _T_2903)) : _T_2903;	// sequencer-master.scala:131:52, :183:52
      wire _T_2912 = io_op_bits_active_vamo ? ~_T_314 & (_T_291 & &_T_0 | _T_2286 & _T_291 | _T_2266 & _T_291 |
                ~_T_291 & ~_T_132 & (_T_2276 & _T_4 | _T_2266 & _T_4 | ~_T_4 & _T_2904)) : _T_2904;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_2913 = io_op_bits_active_vamo ? _T_2308 & _T_314 | ~_T_314 & ~_T_291 & (_T_2308 & _T_132 | ~_T_132
                & ~_T_4 & _T_2881) : _T_2881;	// sequencer-master.scala:132:52, :184:52
      wire _T_2914 = io_op_bits_active_vamo ? _T_2309 & _T_314 | ~_T_314 & ~_T_291 & (_T_2309 & _T_132 | ~_T_132
                & ~_T_4 & _T_2883) : _T_2883;	// sequencer-master.scala:132:52, :184:52
      wire _T_2915 = io_op_bits_active_vamo ? _T_2310 & _T_314 | ~_T_314 & ~_T_291 & (_T_2310 & _T_132 | ~_T_132
                & ~_T_4 & _T_2885) : _T_2885;	// sequencer-master.scala:132:52, :184:52
      wire _T_2916 = io_op_bits_active_vamo ? _T_2311 & _T_314 | ~_T_314 & ~_T_291 & (_T_2311 & _T_132 | ~_T_132
                & ~_T_4 & _T_2887) : _T_2887;	// sequencer-master.scala:132:52, :184:52
      wire _T_2917 = io_op_bits_active_vamo ? _T_2312 & _T_314 | ~_T_314 & ~_T_291 & (_T_2312 & _T_132 | ~_T_132
                & ~_T_4 & _T_2889) : _T_2889;	// sequencer-master.scala:132:52, :184:52
      wire _T_2918 = io_op_bits_active_vamo ? _T_2313 & _T_314 | ~_T_314 & ~_T_291 & (_T_2313 & _T_132 | ~_T_132
                & ~_T_4 & _T_2891) : _T_2891;	// sequencer-master.scala:132:52, :184:52
      wire _T_2919 = io_op_bits_active_vamo ? _T_2314 & _T_314 | ~_T_314 & ~_T_291 & (_T_2314 & _T_132 | ~_T_132
                & ~_T_4 & _T_2893) : _T_2893;	// sequencer-master.scala:132:52, :184:52
      wire _T_2920 = io_op_bits_active_vamo ? _T_2315 & _T_314 | ~_T_314 & ~_T_291 & (_T_2315 & _T_132 | ~_T_132
                & ~_T_4 & _T_2895) : _T_2895;	// sequencer-master.scala:132:52, :184:52
      wire _T_2921 = io_op_bits_active_vamo ? _T_2299 & _T_314 | ~_T_314 & ~_T_291 & (_T_2299 & _T_132 | ~_T_132
                & ~_T_4 & _T_2882) : _T_2882;	// sequencer-master.scala:133:52, :185:52
      wire _T_2922 = io_op_bits_active_vamo ? _T_2300 & _T_314 | ~_T_314 & ~_T_291 & (_T_2300 & _T_132 | ~_T_132
                & ~_T_4 & _T_2884) : _T_2884;	// sequencer-master.scala:133:52, :185:52
      wire _T_2923 = io_op_bits_active_vamo ? _T_2301 & _T_314 | ~_T_314 & ~_T_291 & (_T_2301 & _T_132 | ~_T_132
                & ~_T_4 & _T_2886) : _T_2886;	// sequencer-master.scala:133:52, :185:52
      wire _T_2924 = io_op_bits_active_vamo ? _T_2302 & _T_314 | ~_T_314 & ~_T_291 & (_T_2302 & _T_132 | ~_T_132
                & ~_T_4 & _T_2888) : _T_2888;	// sequencer-master.scala:133:52, :185:52
      wire _T_2925 = io_op_bits_active_vamo ? _T_2303 & _T_314 | ~_T_314 & ~_T_291 & (_T_2303 & _T_132 | ~_T_132
                & ~_T_4 & _T_2890) : _T_2890;	// sequencer-master.scala:133:52, :185:52
      wire _T_2926 = io_op_bits_active_vamo ? _T_2304 & _T_314 | ~_T_314 & ~_T_291 & (_T_2304 & _T_132 | ~_T_132
                & ~_T_4 & _T_2892) : _T_2892;	// sequencer-master.scala:133:52, :185:52
      wire _T_2927 = io_op_bits_active_vamo ? _T_2305 & _T_314 | ~_T_314 & ~_T_291 & (_T_2305 & _T_132 | ~_T_132
                & ~_T_4 & _T_2894) : _T_2894;	// sequencer-master.scala:133:52, :185:52
      wire _T_2928 = io_op_bits_active_vamo ? _T_2306 & _T_314 | ~_T_314 & ~_T_291 & (_T_2306 & _T_132 | ~_T_132
                & ~_T_4 & _T_2896) : _T_2896;	// sequencer-master.scala:133:52, :185:52
      wire _T_2929 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2279 & _T_4 | _T_2238 & _T_4 | ~_T_4 &
                _T_2905) : _T_2905;	// sequencer-master.scala:131:52, :183:52
      wire _T_2930 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2280 & _T_4 | _T_2242 & _T_4 | ~_T_4 &
                _T_2906) : _T_2906;	// sequencer-master.scala:131:52, :183:52
      wire _T_2931 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2281 & _T_4 | _T_2246 & _T_4 | ~_T_4 &
                _T_2907) : _T_2907;	// sequencer-master.scala:131:52, :183:52
      wire _T_2932 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2282 & _T_4 | _T_2250 & _T_4 | ~_T_4 &
                _T_2908) : _T_2908;	// sequencer-master.scala:131:52, :183:52
      wire _T_2933 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2283 & _T_4 | _T_2254 & _T_4 | ~_T_4 &
                _T_2909) : _T_2909;	// sequencer-master.scala:131:52, :183:52
      wire _T_2934 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2284 & _T_4 | _T_2258 & _T_4 | ~_T_4 &
                _T_2910) : _T_2910;	// sequencer-master.scala:131:52, :183:52
      wire _T_2935 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2285 & _T_4 | _T_2262 & _T_4 | ~_T_4 &
                _T_2911) : _T_2911;	// sequencer-master.scala:131:52, :183:52
      wire _T_2936 = io_op_bits_active_vldx ? ~_T_291 & ~_T_132 & (_T_2286 & _T_4 | _T_2266 & _T_4 | ~_T_4 &
                _T_2912) : _T_2912;	// sequencer-master.scala:131:52, :183:52
      wire _T_2937 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2308 &
                _T_291 | ~_T_291 & (_T_2308 & _T_132 | ~_T_132 & ~_T_4 & _T_2913) : _T_2913);	// sequencer-master.scala:132:52, :184:52
      wire _T_2938 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2299 &
                _T_291 | ~_T_291 & (_T_2299 & _T_132 | ~_T_132 & ~_T_4 & _T_2921) : _T_2921);	// sequencer-master.scala:133:52, :185:52
      wire _T_2939 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2309 &
                _T_291 | ~_T_291 & (_T_2309 & _T_132 | ~_T_132 & ~_T_4 & _T_2914) : _T_2914);	// sequencer-master.scala:132:52, :184:52
      wire _T_2940 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2300 &
                _T_291 | ~_T_291 & (_T_2300 & _T_132 | ~_T_132 & ~_T_4 & _T_2922) : _T_2922);	// sequencer-master.scala:133:52, :185:52
      wire _T_2941 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2310 &
                _T_291 | ~_T_291 & (_T_2310 & _T_132 | ~_T_132 & ~_T_4 & _T_2915) : _T_2915);	// sequencer-master.scala:132:52, :184:52
      wire _T_2942 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2301 &
                _T_291 | ~_T_291 & (_T_2301 & _T_132 | ~_T_132 & ~_T_4 & _T_2923) : _T_2923);	// sequencer-master.scala:133:52, :185:52
      wire _T_2943 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2311 &
                _T_291 | ~_T_291 & (_T_2311 & _T_132 | ~_T_132 & ~_T_4 & _T_2916) : _T_2916);	// sequencer-master.scala:132:52, :184:52
      wire _T_2944 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2302 &
                _T_291 | ~_T_291 & (_T_2302 & _T_132 | ~_T_132 & ~_T_4 & _T_2924) : _T_2924);	// sequencer-master.scala:133:52, :185:52
      wire _T_2945 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2312 &
                _T_291 | ~_T_291 & (_T_2312 & _T_132 | ~_T_132 & ~_T_4 & _T_2917) : _T_2917);	// sequencer-master.scala:132:52, :184:52
      wire _T_2946 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2303 &
                _T_291 | ~_T_291 & (_T_2303 & _T_132 | ~_T_132 & ~_T_4 & _T_2925) : _T_2925);	// sequencer-master.scala:133:52, :185:52
      wire _T_2947 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2313 &
                _T_291 | ~_T_291 & (_T_2313 & _T_132 | ~_T_132 & ~_T_4 & _T_2918) : _T_2918);	// sequencer-master.scala:132:52, :184:52
      wire _T_2948 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2304 &
                _T_291 | ~_T_291 & (_T_2304 & _T_132 | ~_T_132 & ~_T_4 & _T_2926) : _T_2926);	// sequencer-master.scala:133:52, :185:52
      wire _T_2949 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2314 &
                _T_291 | ~_T_291 & (_T_2314 & _T_132 | ~_T_132 & ~_T_4 & _T_2919) : _T_2919);	// sequencer-master.scala:132:52, :184:52
      wire _T_2950 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2305 &
                _T_291 | ~_T_291 & (_T_2305 & _T_132 | ~_T_132 & ~_T_4 & _T_2927) : _T_2927);	// sequencer-master.scala:133:52, :185:52
      wire _T_2951 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2315 &
                _T_291 | ~_T_291 & (_T_2315 & _T_132 | ~_T_132 & ~_T_4 & _T_2920) : _T_2920);	// sequencer-master.scala:132:52, :184:52
      wire _T_2952 = (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vldx ? _T_2306 &
                _T_291 | ~_T_291 & (_T_2306 & _T_132 | ~_T_132 & ~_T_4 & _T_2928) : _T_2928);	// sequencer-master.scala:133:52, :185:52
      wire _T_2953 = io_op_bits_active_vstx ? _T_291 & _T_132 | _T_2299 & _T_291 | _T_2238 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2279 & _T_4 | _T_2238 & _T_4 | ~_T_4 & _T_2929) : _T_2929;	// sequencer-master.scala:131:52, :183:52
      wire _T_2954 = io_op_bits_active_vstx ? _T_291 & _T_133 | _T_2300 & _T_291 | _T_2242 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2280 & _T_4 | _T_2242 & _T_4 | ~_T_4 & _T_2930) : _T_2930;	// sequencer-master.scala:131:52, :183:52
      wire _T_2955 = io_op_bits_active_vstx ? _T_291 & _T_134 | _T_2301 & _T_291 | _T_2246 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2281 & _T_4 | _T_2246 & _T_4 | ~_T_4 & _T_2931) : _T_2931;	// sequencer-master.scala:131:52, :183:52
      wire _T_2956 = io_op_bits_active_vstx ? _T_291 & _T_135 | _T_2302 & _T_291 | _T_2250 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2282 & _T_4 | _T_2250 & _T_4 | ~_T_4 & _T_2932) : _T_2932;	// sequencer-master.scala:131:52, :183:52
      wire _T_2957 = io_op_bits_active_vstx ? _T_291 & _T_136 | _T_2303 & _T_291 | _T_2254 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2283 & _T_4 | _T_2254 & _T_4 | ~_T_4 & _T_2933) : _T_2933;	// sequencer-master.scala:131:52, :183:52
      wire _T_2958 = io_op_bits_active_vstx ? _T_291 & _T_137 | _T_2304 & _T_291 | _T_2258 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2284 & _T_4 | _T_2258 & _T_4 | ~_T_4 & _T_2934) : _T_2934;	// sequencer-master.scala:131:52, :183:52
      wire _T_2959 = io_op_bits_active_vstx ? _T_291 & _T_138 | _T_2305 & _T_291 | _T_2262 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2285 & _T_4 | _T_2262 & _T_4 | ~_T_4 & _T_2935) : _T_2935;	// sequencer-master.scala:131:52, :183:52
      wire _T_2960 = io_op_bits_active_vstx ? _T_291 & &_T_0 | _T_2306 & _T_291 | _T_2266 & _T_291 | ~_T_291 &
                ~_T_132 & (_T_2286 & _T_4 | _T_2266 & _T_4 | ~_T_4 & _T_2936) : _T_2936;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_2961 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2238 & _T_4 | ~_T_4 & _T_2953) : _T_2953;	// sequencer-master.scala:131:52, :183:52
      wire _T_2962 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2242 & _T_4 | ~_T_4 & _T_2954) : _T_2954;	// sequencer-master.scala:131:52, :183:52
      wire _T_2963 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2246 & _T_4 | ~_T_4 & _T_2955) : _T_2955;	// sequencer-master.scala:131:52, :183:52
      wire _T_2964 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2250 & _T_4 | ~_T_4 & _T_2956) : _T_2956;	// sequencer-master.scala:131:52, :183:52
      wire _T_2965 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2254 & _T_4 | ~_T_4 & _T_2957) : _T_2957;	// sequencer-master.scala:131:52, :183:52
      wire _T_2966 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2258 & _T_4 | ~_T_4 & _T_2958) : _T_2958;	// sequencer-master.scala:131:52, :183:52
      wire _T_2967 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2262 & _T_4 | ~_T_4 & _T_2959) : _T_2959;	// sequencer-master.scala:131:52, :183:52
      wire _T_2968 = io_op_bits_active_vld ? ~_T_291 & ~_T_132 & (_T_2266 & _T_4 | ~_T_4 & _T_2960) : _T_2960;	// sequencer-master.scala:131:52, :183:52
      wire _T_2969 = io_op_bits_active_vint ? _T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 &
                e_1_raw_0 : e_1_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_2970 = io_op_bits_active_vint ? _T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 &
                e_1_raw_1 : e_1_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_2971 = io_op_bits_active_vint ? _T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 &
                e_1_raw_2 : e_1_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_2972 = io_op_bits_active_vint ? _T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 &
                e_1_raw_3 : e_1_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_2973 = io_op_bits_active_vint ? _T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 &
                e_1_raw_4 : e_1_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_2974 = io_op_bits_active_vint ? _T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 &
                e_1_raw_5 : e_1_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_2975 = io_op_bits_active_vint ? _T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 &
                e_1_raw_6 : e_1_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_2976 = io_op_bits_active_vint ? _T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 &
                e_1_raw_7 : e_1_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_2977 = io_op_bits_active_vint ? _T_2308 & _T_5 | ~_T_5 & e_1_war_0 : e_1_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_2978 = io_op_bits_active_vint ? _T_2309 & _T_5 | ~_T_5 & e_1_war_1 : e_1_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_2979 = io_op_bits_active_vint ? _T_2310 & _T_5 | ~_T_5 & e_1_war_2 : e_1_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_2980 = io_op_bits_active_vint ? _T_2311 & _T_5 | ~_T_5 & e_1_war_3 : e_1_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_2981 = io_op_bits_active_vint ? _T_2312 & _T_5 | ~_T_5 & e_1_war_4 : e_1_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_2982 = io_op_bits_active_vint ? _T_2313 & _T_5 | ~_T_5 & e_1_war_5 : e_1_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_2983 = io_op_bits_active_vint ? _T_2314 & _T_5 | ~_T_5 & e_1_war_6 : e_1_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_2984 = io_op_bits_active_vint ? _T_2315 & _T_5 | ~_T_5 & e_1_war_7 : e_1_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_2985 = io_op_bits_active_vint ? _T_2299 & _T_5 | ~_T_5 & e_1_waw_0 : e_1_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_2986 = io_op_bits_active_vint ? _T_2300 & _T_5 | ~_T_5 & e_1_waw_1 : e_1_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_2987 = io_op_bits_active_vint ? _T_2301 & _T_5 | ~_T_5 & e_1_waw_2 : e_1_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_2988 = io_op_bits_active_vint ? _T_2302 & _T_5 | ~_T_5 & e_1_waw_3 : e_1_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_2989 = io_op_bits_active_vint ? _T_2303 & _T_5 | ~_T_5 & e_1_waw_4 : e_1_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_2990 = io_op_bits_active_vint ? _T_2304 & _T_5 | ~_T_5 & e_1_waw_5 : e_1_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_2991 = io_op_bits_active_vint ? _T_2305 & _T_5 | ~_T_5 & e_1_waw_6 : e_1_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_2992 = io_op_bits_active_vint ? _T_2306 & _T_5 | ~_T_5 & e_1_waw_7 : e_1_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_2993 = io_op_bits_active_vipred ? _T_2289 & _T_5 | _T_2279 & _T_5 | _T_2269 & _T_5 | ~_T_5 &
                _T_2969 : _T_2969;	// sequencer-master.scala:131:52, :183:52
      wire _T_2994 = io_op_bits_active_vipred ? _T_2290 & _T_5 | _T_2280 & _T_5 | _T_2270 & _T_5 | ~_T_5 &
                _T_2970 : _T_2970;	// sequencer-master.scala:131:52, :183:52
      wire _T_2995 = io_op_bits_active_vipred ? _T_2291 & _T_5 | _T_2281 & _T_5 | _T_2271 & _T_5 | ~_T_5 &
                _T_2971 : _T_2971;	// sequencer-master.scala:131:52, :183:52
      wire _T_2996 = io_op_bits_active_vipred ? _T_2292 & _T_5 | _T_2282 & _T_5 | _T_2272 & _T_5 | ~_T_5 &
                _T_2972 : _T_2972;	// sequencer-master.scala:131:52, :183:52
      wire _T_2997 = io_op_bits_active_vipred ? _T_2293 & _T_5 | _T_2283 & _T_5 | _T_2273 & _T_5 | ~_T_5 &
                _T_2973 : _T_2973;	// sequencer-master.scala:131:52, :183:52
      wire _T_2998 = io_op_bits_active_vipred ? _T_2294 & _T_5 | _T_2284 & _T_5 | _T_2274 & _T_5 | ~_T_5 &
                _T_2974 : _T_2974;	// sequencer-master.scala:131:52, :183:52
      wire _T_2999 = io_op_bits_active_vipred ? _T_2295 & _T_5 | _T_2285 & _T_5 | _T_2275 & _T_5 | ~_T_5 &
                _T_2975 : _T_2975;	// sequencer-master.scala:131:52, :183:52
      wire _T_3000 = io_op_bits_active_vipred ? _T_2296 & _T_5 | _T_2286 & _T_5 | _T_2276 & _T_5 | ~_T_5 &
                _T_2976 : _T_2976;	// sequencer-master.scala:131:52, :183:52
      wire _T_3001 = io_op_bits_active_vipred ? _T_2308 & _T_5 | ~_T_5 & _T_2977 : _T_2977;	// sequencer-master.scala:132:52, :184:52
      wire _T_3002 = io_op_bits_active_vipred ? _T_2309 & _T_5 | ~_T_5 & _T_2978 : _T_2978;	// sequencer-master.scala:132:52, :184:52
      wire _T_3003 = io_op_bits_active_vipred ? _T_2310 & _T_5 | ~_T_5 & _T_2979 : _T_2979;	// sequencer-master.scala:132:52, :184:52
      wire _T_3004 = io_op_bits_active_vipred ? _T_2311 & _T_5 | ~_T_5 & _T_2980 : _T_2980;	// sequencer-master.scala:132:52, :184:52
      wire _T_3005 = io_op_bits_active_vipred ? _T_2312 & _T_5 | ~_T_5 & _T_2981 : _T_2981;	// sequencer-master.scala:132:52, :184:52
      wire _T_3006 = io_op_bits_active_vipred ? _T_2313 & _T_5 | ~_T_5 & _T_2982 : _T_2982;	// sequencer-master.scala:132:52, :184:52
      wire _T_3007 = io_op_bits_active_vipred ? _T_2314 & _T_5 | ~_T_5 & _T_2983 : _T_2983;	// sequencer-master.scala:132:52, :184:52
      wire _T_3008 = io_op_bits_active_vipred ? _T_2315 & _T_5 | ~_T_5 & _T_2984 : _T_2984;	// sequencer-master.scala:132:52, :184:52
      wire _T_3009 = io_op_bits_active_vipred ? _T_2299 & _T_5 | ~_T_5 & _T_2985 : _T_2985;	// sequencer-master.scala:133:52, :185:52
      wire _T_3010 = io_op_bits_active_vipred ? _T_2300 & _T_5 | ~_T_5 & _T_2986 : _T_2986;	// sequencer-master.scala:133:52, :185:52
      wire _T_3011 = io_op_bits_active_vipred ? _T_2301 & _T_5 | ~_T_5 & _T_2987 : _T_2987;	// sequencer-master.scala:133:52, :185:52
      wire _T_3012 = io_op_bits_active_vipred ? _T_2302 & _T_5 | ~_T_5 & _T_2988 : _T_2988;	// sequencer-master.scala:133:52, :185:52
      wire _T_3013 = io_op_bits_active_vipred ? _T_2303 & _T_5 | ~_T_5 & _T_2989 : _T_2989;	// sequencer-master.scala:133:52, :185:52
      wire _T_3014 = io_op_bits_active_vipred ? _T_2304 & _T_5 | ~_T_5 & _T_2990 : _T_2990;	// sequencer-master.scala:133:52, :185:52
      wire _T_3015 = io_op_bits_active_vipred ? _T_2305 & _T_5 | ~_T_5 & _T_2991 : _T_2991;	// sequencer-master.scala:133:52, :185:52
      wire _T_3016 = io_op_bits_active_vipred ? _T_2306 & _T_5 | ~_T_5 & _T_2992 : _T_2992;	// sequencer-master.scala:133:52, :185:52
      wire _T_3017 = io_op_bits_active_vimul ? _T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 &
                _T_2993 : _T_2993;	// sequencer-master.scala:131:52, :183:52
      wire _T_3018 = io_op_bits_active_vimul ? _T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 &
                _T_2994 : _T_2994;	// sequencer-master.scala:131:52, :183:52
      wire _T_3019 = io_op_bits_active_vimul ? _T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 &
                _T_2995 : _T_2995;	// sequencer-master.scala:131:52, :183:52
      wire _T_3020 = io_op_bits_active_vimul ? _T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 &
                _T_2996 : _T_2996;	// sequencer-master.scala:131:52, :183:52
      wire _T_3021 = io_op_bits_active_vimul ? _T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 &
                _T_2997 : _T_2997;	// sequencer-master.scala:131:52, :183:52
      wire _T_3022 = io_op_bits_active_vimul ? _T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 &
                _T_2998 : _T_2998;	// sequencer-master.scala:131:52, :183:52
      wire _T_3023 = io_op_bits_active_vimul ? _T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 &
                _T_2999 : _T_2999;	// sequencer-master.scala:131:52, :183:52
      wire _T_3024 = io_op_bits_active_vimul ? _T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 &
                _T_3000 : _T_3000;	// sequencer-master.scala:131:52, :183:52
      wire _T_3025 = io_op_bits_active_vimul ? _T_2308 & _T_5 | ~_T_5 & _T_3001 : _T_3001;	// sequencer-master.scala:132:52, :184:52
      wire _T_3026 = io_op_bits_active_vimul ? _T_2309 & _T_5 | ~_T_5 & _T_3002 : _T_3002;	// sequencer-master.scala:132:52, :184:52
      wire _T_3027 = io_op_bits_active_vimul ? _T_2310 & _T_5 | ~_T_5 & _T_3003 : _T_3003;	// sequencer-master.scala:132:52, :184:52
      wire _T_3028 = io_op_bits_active_vimul ? _T_2311 & _T_5 | ~_T_5 & _T_3004 : _T_3004;	// sequencer-master.scala:132:52, :184:52
      wire _T_3029 = io_op_bits_active_vimul ? _T_2312 & _T_5 | ~_T_5 & _T_3005 : _T_3005;	// sequencer-master.scala:132:52, :184:52
      wire _T_3030 = io_op_bits_active_vimul ? _T_2313 & _T_5 | ~_T_5 & _T_3006 : _T_3006;	// sequencer-master.scala:132:52, :184:52
      wire _T_3031 = io_op_bits_active_vimul ? _T_2314 & _T_5 | ~_T_5 & _T_3007 : _T_3007;	// sequencer-master.scala:132:52, :184:52
      wire _T_3032 = io_op_bits_active_vimul ? _T_2315 & _T_5 | ~_T_5 & _T_3008 : _T_3008;	// sequencer-master.scala:132:52, :184:52
      wire _T_3033 = io_op_bits_active_vimul ? _T_2299 & _T_5 | ~_T_5 & _T_3009 : _T_3009;	// sequencer-master.scala:133:52, :185:52
      wire _T_3034 = io_op_bits_active_vimul ? _T_2300 & _T_5 | ~_T_5 & _T_3010 : _T_3010;	// sequencer-master.scala:133:52, :185:52
      wire _T_3035 = io_op_bits_active_vimul ? _T_2301 & _T_5 | ~_T_5 & _T_3011 : _T_3011;	// sequencer-master.scala:133:52, :185:52
      wire _T_3036 = io_op_bits_active_vimul ? _T_2302 & _T_5 | ~_T_5 & _T_3012 : _T_3012;	// sequencer-master.scala:133:52, :185:52
      wire _T_3037 = io_op_bits_active_vimul ? _T_2303 & _T_5 | ~_T_5 & _T_3013 : _T_3013;	// sequencer-master.scala:133:52, :185:52
      wire _T_3038 = io_op_bits_active_vimul ? _T_2304 & _T_5 | ~_T_5 & _T_3014 : _T_3014;	// sequencer-master.scala:133:52, :185:52
      wire _T_3039 = io_op_bits_active_vimul ? _T_2305 & _T_5 | ~_T_5 & _T_3015 : _T_3015;	// sequencer-master.scala:133:52, :185:52
      wire _T_3040 = io_op_bits_active_vimul ? _T_2306 & _T_5 | ~_T_5 & _T_3016 : _T_3016;	// sequencer-master.scala:133:52, :185:52
      wire _T_3041 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5 |
                ~_T_5 & _T_3017) : _T_3017;	// sequencer-master.scala:131:52, :183:52
      wire _T_3042 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5 |
                ~_T_5 & _T_3018) : _T_3018;	// sequencer-master.scala:131:52, :183:52
      wire _T_3043 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5 |
                ~_T_5 & _T_3019) : _T_3019;	// sequencer-master.scala:131:52, :183:52
      wire _T_3044 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5 |
                ~_T_5 & _T_3020) : _T_3020;	// sequencer-master.scala:131:52, :183:52
      wire _T_3045 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5 |
                ~_T_5 & _T_3021) : _T_3021;	// sequencer-master.scala:131:52, :183:52
      wire _T_3046 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5 |
                ~_T_5 & _T_3022) : _T_3022;	// sequencer-master.scala:131:52, :183:52
      wire _T_3047 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5 |
                ~_T_5 & _T_3023) : _T_3023;	// sequencer-master.scala:131:52, :183:52
      wire _T_3048 = io_op_bits_active_vidiv ? ~_T_133 & (_T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5 |
                ~_T_5 & _T_3024) : _T_3024;	// sequencer-master.scala:131:52, :183:52
      wire _T_3049 = io_op_bits_active_vidiv ? _T_2308 & _T_133 | ~_T_133 & (_T_2308 & _T_5 | ~_T_5 & _T_3025) :
                _T_3025;	// sequencer-master.scala:132:52, :184:52
      wire _T_3050 = io_op_bits_active_vidiv ? _T_2309 & _T_133 | ~_T_133 & (_T_2309 & _T_5 | ~_T_5 & _T_3026) :
                _T_3026;	// sequencer-master.scala:132:52, :184:52
      wire _T_3051 = io_op_bits_active_vidiv ? _T_2310 & _T_133 | ~_T_133 & (_T_2310 & _T_5 | ~_T_5 & _T_3027) :
                _T_3027;	// sequencer-master.scala:132:52, :184:52
      wire _T_3052 = io_op_bits_active_vidiv ? _T_2311 & _T_133 | ~_T_133 & (_T_2311 & _T_5 | ~_T_5 & _T_3028) :
                _T_3028;	// sequencer-master.scala:132:52, :184:52
      wire _T_3053 = io_op_bits_active_vidiv ? _T_2312 & _T_133 | ~_T_133 & (_T_2312 & _T_5 | ~_T_5 & _T_3029) :
                _T_3029;	// sequencer-master.scala:132:52, :184:52
      wire _T_3054 = io_op_bits_active_vidiv ? _T_2313 & _T_133 | ~_T_133 & (_T_2313 & _T_5 | ~_T_5 & _T_3030) :
                _T_3030;	// sequencer-master.scala:132:52, :184:52
      wire _T_3055 = io_op_bits_active_vidiv ? _T_2314 & _T_133 | ~_T_133 & (_T_2314 & _T_5 | ~_T_5 & _T_3031) :
                _T_3031;	// sequencer-master.scala:132:52, :184:52
      wire _T_3056 = io_op_bits_active_vidiv ? _T_2315 & _T_133 | ~_T_133 & (_T_2315 & _T_5 | ~_T_5 & _T_3032) :
                _T_3032;	// sequencer-master.scala:132:52, :184:52
      wire _T_3057 = io_op_bits_active_vidiv ? _T_2299 & _T_133 | ~_T_133 & (_T_2299 & _T_5 | ~_T_5 & _T_3033) :
                _T_3033;	// sequencer-master.scala:133:52, :185:52
      wire _T_3058 = io_op_bits_active_vidiv ? _T_2300 & _T_133 | ~_T_133 & (_T_2300 & _T_5 | ~_T_5 & _T_3034) :
                _T_3034;	// sequencer-master.scala:133:52, :185:52
      wire _T_3059 = io_op_bits_active_vidiv ? _T_2301 & _T_133 | ~_T_133 & (_T_2301 & _T_5 | ~_T_5 & _T_3035) :
                _T_3035;	// sequencer-master.scala:133:52, :185:52
      wire _T_3060 = io_op_bits_active_vidiv ? _T_2302 & _T_133 | ~_T_133 & (_T_2302 & _T_5 | ~_T_5 & _T_3036) :
                _T_3036;	// sequencer-master.scala:133:52, :185:52
      wire _T_3061 = io_op_bits_active_vidiv ? _T_2303 & _T_133 | ~_T_133 & (_T_2303 & _T_5 | ~_T_5 & _T_3037) :
                _T_3037;	// sequencer-master.scala:133:52, :185:52
      wire _T_3062 = io_op_bits_active_vidiv ? _T_2304 & _T_133 | ~_T_133 & (_T_2304 & _T_5 | ~_T_5 & _T_3038) :
                _T_3038;	// sequencer-master.scala:133:52, :185:52
      wire _T_3063 = io_op_bits_active_vidiv ? _T_2305 & _T_133 | ~_T_133 & (_T_2305 & _T_5 | ~_T_5 & _T_3039) :
                _T_3039;	// sequencer-master.scala:133:52, :185:52
      wire _T_3064 = io_op_bits_active_vidiv ? _T_2306 & _T_133 | ~_T_133 & (_T_2306 & _T_5 | ~_T_5 & _T_3040) :
                _T_3040;	// sequencer-master.scala:133:52, :185:52
      wire _T_3065 = io_op_bits_active_vfma ? _T_2289 & _T_5 | _T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5
                | ~_T_5 & _T_3041 : _T_3041;	// sequencer-master.scala:131:52, :183:52
      wire _T_3066 = io_op_bits_active_vfma ? _T_2290 & _T_5 | _T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5
                | ~_T_5 & _T_3042 : _T_3042;	// sequencer-master.scala:131:52, :183:52
      wire _T_3067 = io_op_bits_active_vfma ? _T_2291 & _T_5 | _T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5
                | ~_T_5 & _T_3043 : _T_3043;	// sequencer-master.scala:131:52, :183:52
      wire _T_3068 = io_op_bits_active_vfma ? _T_2292 & _T_5 | _T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5
                | ~_T_5 & _T_3044 : _T_3044;	// sequencer-master.scala:131:52, :183:52
      wire _T_3069 = io_op_bits_active_vfma ? _T_2293 & _T_5 | _T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5
                | ~_T_5 & _T_3045 : _T_3045;	// sequencer-master.scala:131:52, :183:52
      wire _T_3070 = io_op_bits_active_vfma ? _T_2294 & _T_5 | _T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5
                | ~_T_5 & _T_3046 : _T_3046;	// sequencer-master.scala:131:52, :183:52
      wire _T_3071 = io_op_bits_active_vfma ? _T_2295 & _T_5 | _T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5
                | ~_T_5 & _T_3047 : _T_3047;	// sequencer-master.scala:131:52, :183:52
      wire _T_3072 = io_op_bits_active_vfma ? _T_2296 & _T_5 | _T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5
                | ~_T_5 & _T_3048 : _T_3048;	// sequencer-master.scala:131:52, :183:52
      wire _T_3073 = io_op_bits_active_vfma ? _T_2308 & _T_5 | ~_T_5 & _T_3049 : _T_3049;	// sequencer-master.scala:132:52, :184:52
      wire _T_3074 = io_op_bits_active_vfma ? _T_2309 & _T_5 | ~_T_5 & _T_3050 : _T_3050;	// sequencer-master.scala:132:52, :184:52
      wire _T_3075 = io_op_bits_active_vfma ? _T_2310 & _T_5 | ~_T_5 & _T_3051 : _T_3051;	// sequencer-master.scala:132:52, :184:52
      wire _T_3076 = io_op_bits_active_vfma ? _T_2311 & _T_5 | ~_T_5 & _T_3052 : _T_3052;	// sequencer-master.scala:132:52, :184:52
      wire _T_3077 = io_op_bits_active_vfma ? _T_2312 & _T_5 | ~_T_5 & _T_3053 : _T_3053;	// sequencer-master.scala:132:52, :184:52
      wire _T_3078 = io_op_bits_active_vfma ? _T_2313 & _T_5 | ~_T_5 & _T_3054 : _T_3054;	// sequencer-master.scala:132:52, :184:52
      wire _T_3079 = io_op_bits_active_vfma ? _T_2314 & _T_5 | ~_T_5 & _T_3055 : _T_3055;	// sequencer-master.scala:132:52, :184:52
      wire _T_3080 = io_op_bits_active_vfma ? _T_2315 & _T_5 | ~_T_5 & _T_3056 : _T_3056;	// sequencer-master.scala:132:52, :184:52
      wire _T_3081 = io_op_bits_active_vfma ? _T_2299 & _T_5 | ~_T_5 & _T_3057 : _T_3057;	// sequencer-master.scala:133:52, :185:52
      wire _T_3082 = io_op_bits_active_vfma ? _T_2300 & _T_5 | ~_T_5 & _T_3058 : _T_3058;	// sequencer-master.scala:133:52, :185:52
      wire _T_3083 = io_op_bits_active_vfma ? _T_2301 & _T_5 | ~_T_5 & _T_3059 : _T_3059;	// sequencer-master.scala:133:52, :185:52
      wire _T_3084 = io_op_bits_active_vfma ? _T_2302 & _T_5 | ~_T_5 & _T_3060 : _T_3060;	// sequencer-master.scala:133:52, :185:52
      wire _T_3085 = io_op_bits_active_vfma ? _T_2303 & _T_5 | ~_T_5 & _T_3061 : _T_3061;	// sequencer-master.scala:133:52, :185:52
      wire _T_3086 = io_op_bits_active_vfma ? _T_2304 & _T_5 | ~_T_5 & _T_3062 : _T_3062;	// sequencer-master.scala:133:52, :185:52
      wire _T_3087 = io_op_bits_active_vfma ? _T_2305 & _T_5 | ~_T_5 & _T_3063 : _T_3063;	// sequencer-master.scala:133:52, :185:52
      wire _T_3088 = io_op_bits_active_vfma ? _T_2306 & _T_5 | ~_T_5 & _T_3064 : _T_3064;	// sequencer-master.scala:133:52, :185:52
      wire _T_3089 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5 |
                ~_T_5 & _T_3065) : _T_3065;	// sequencer-master.scala:131:52, :183:52
      wire _T_3090 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5 |
                ~_T_5 & _T_3066) : _T_3066;	// sequencer-master.scala:131:52, :183:52
      wire _T_3091 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5 |
                ~_T_5 & _T_3067) : _T_3067;	// sequencer-master.scala:131:52, :183:52
      wire _T_3092 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5 |
                ~_T_5 & _T_3068) : _T_3068;	// sequencer-master.scala:131:52, :183:52
      wire _T_3093 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5 |
                ~_T_5 & _T_3069) : _T_3069;	// sequencer-master.scala:131:52, :183:52
      wire _T_3094 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5 |
                ~_T_5 & _T_3070) : _T_3070;	// sequencer-master.scala:131:52, :183:52
      wire _T_3095 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5 |
                ~_T_5 & _T_3071) : _T_3071;	// sequencer-master.scala:131:52, :183:52
      wire _T_3096 = io_op_bits_active_vfdiv ? ~_T_133 & (_T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5 |
                ~_T_5 & _T_3072) : _T_3072;	// sequencer-master.scala:131:52, :183:52
      wire _T_3097 = io_op_bits_active_vfdiv ? _T_2308 & _T_133 | ~_T_133 & (_T_2308 & _T_5 | ~_T_5 & _T_3073) :
                _T_3073;	// sequencer-master.scala:132:52, :184:52
      wire _T_3098 = io_op_bits_active_vfdiv ? _T_2309 & _T_133 | ~_T_133 & (_T_2309 & _T_5 | ~_T_5 & _T_3074) :
                _T_3074;	// sequencer-master.scala:132:52, :184:52
      wire _T_3099 = io_op_bits_active_vfdiv ? _T_2310 & _T_133 | ~_T_133 & (_T_2310 & _T_5 | ~_T_5 & _T_3075) :
                _T_3075;	// sequencer-master.scala:132:52, :184:52
      wire _T_3100 = io_op_bits_active_vfdiv ? _T_2311 & _T_133 | ~_T_133 & (_T_2311 & _T_5 | ~_T_5 & _T_3076) :
                _T_3076;	// sequencer-master.scala:132:52, :184:52
      wire _T_3101 = io_op_bits_active_vfdiv ? _T_2312 & _T_133 | ~_T_133 & (_T_2312 & _T_5 | ~_T_5 & _T_3077) :
                _T_3077;	// sequencer-master.scala:132:52, :184:52
      wire _T_3102 = io_op_bits_active_vfdiv ? _T_2313 & _T_133 | ~_T_133 & (_T_2313 & _T_5 | ~_T_5 & _T_3078) :
                _T_3078;	// sequencer-master.scala:132:52, :184:52
      wire _T_3103 = io_op_bits_active_vfdiv ? _T_2314 & _T_133 | ~_T_133 & (_T_2314 & _T_5 | ~_T_5 & _T_3079) :
                _T_3079;	// sequencer-master.scala:132:52, :184:52
      wire _T_3104 = io_op_bits_active_vfdiv ? _T_2315 & _T_133 | ~_T_133 & (_T_2315 & _T_5 | ~_T_5 & _T_3080) :
                _T_3080;	// sequencer-master.scala:132:52, :184:52
      wire _T_3105 = io_op_bits_active_vfdiv ? _T_2299 & _T_133 | ~_T_133 & (_T_2299 & _T_5 | ~_T_5 & _T_3081) :
                _T_3081;	// sequencer-master.scala:133:52, :185:52
      wire _T_3106 = io_op_bits_active_vfdiv ? _T_2300 & _T_133 | ~_T_133 & (_T_2300 & _T_5 | ~_T_5 & _T_3082) :
                _T_3082;	// sequencer-master.scala:133:52, :185:52
      wire _T_3107 = io_op_bits_active_vfdiv ? _T_2301 & _T_133 | ~_T_133 & (_T_2301 & _T_5 | ~_T_5 & _T_3083) :
                _T_3083;	// sequencer-master.scala:133:52, :185:52
      wire _T_3108 = io_op_bits_active_vfdiv ? _T_2302 & _T_133 | ~_T_133 & (_T_2302 & _T_5 | ~_T_5 & _T_3084) :
                _T_3084;	// sequencer-master.scala:133:52, :185:52
      wire _T_3109 = io_op_bits_active_vfdiv ? _T_2303 & _T_133 | ~_T_133 & (_T_2303 & _T_5 | ~_T_5 & _T_3085) :
                _T_3085;	// sequencer-master.scala:133:52, :185:52
      wire _T_3110 = io_op_bits_active_vfdiv ? _T_2304 & _T_133 | ~_T_133 & (_T_2304 & _T_5 | ~_T_5 & _T_3086) :
                _T_3086;	// sequencer-master.scala:133:52, :185:52
      wire _T_3111 = io_op_bits_active_vfdiv ? _T_2305 & _T_133 | ~_T_133 & (_T_2305 & _T_5 | ~_T_5 & _T_3087) :
                _T_3087;	// sequencer-master.scala:133:52, :185:52
      wire _T_3112 = io_op_bits_active_vfdiv ? _T_2306 & _T_133 | ~_T_133 & (_T_2306 & _T_5 | ~_T_5 & _T_3088) :
                _T_3088;	// sequencer-master.scala:133:52, :185:52
      wire _T_3113 = io_op_bits_active_vfcmp ? _T_2279 & _T_5 | _T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 &
                _T_3089 : _T_3089;	// sequencer-master.scala:131:52, :183:52
      wire _T_3114 = io_op_bits_active_vfcmp ? _T_2280 & _T_5 | _T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 &
                _T_3090 : _T_3090;	// sequencer-master.scala:131:52, :183:52
      wire _T_3115 = io_op_bits_active_vfcmp ? _T_2281 & _T_5 | _T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 &
                _T_3091 : _T_3091;	// sequencer-master.scala:131:52, :183:52
      wire _T_3116 = io_op_bits_active_vfcmp ? _T_2282 & _T_5 | _T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 &
                _T_3092 : _T_3092;	// sequencer-master.scala:131:52, :183:52
      wire _T_3117 = io_op_bits_active_vfcmp ? _T_2283 & _T_5 | _T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 &
                _T_3093 : _T_3093;	// sequencer-master.scala:131:52, :183:52
      wire _T_3118 = io_op_bits_active_vfcmp ? _T_2284 & _T_5 | _T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 &
                _T_3094 : _T_3094;	// sequencer-master.scala:131:52, :183:52
      wire _T_3119 = io_op_bits_active_vfcmp ? _T_2285 & _T_5 | _T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 &
                _T_3095 : _T_3095;	// sequencer-master.scala:131:52, :183:52
      wire _T_3120 = io_op_bits_active_vfcmp ? _T_2286 & _T_5 | _T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 &
                _T_3096 : _T_3096;	// sequencer-master.scala:131:52, :183:52
      wire _T_3121 = io_op_bits_active_vfcmp ? _T_2308 & _T_5 | ~_T_5 & _T_3097 : _T_3097;	// sequencer-master.scala:132:52, :184:52
      wire _T_3122 = io_op_bits_active_vfcmp ? _T_2309 & _T_5 | ~_T_5 & _T_3098 : _T_3098;	// sequencer-master.scala:132:52, :184:52
      wire _T_3123 = io_op_bits_active_vfcmp ? _T_2310 & _T_5 | ~_T_5 & _T_3099 : _T_3099;	// sequencer-master.scala:132:52, :184:52
      wire _T_3124 = io_op_bits_active_vfcmp ? _T_2311 & _T_5 | ~_T_5 & _T_3100 : _T_3100;	// sequencer-master.scala:132:52, :184:52
      wire _T_3125 = io_op_bits_active_vfcmp ? _T_2312 & _T_5 | ~_T_5 & _T_3101 : _T_3101;	// sequencer-master.scala:132:52, :184:52
      wire _T_3126 = io_op_bits_active_vfcmp ? _T_2313 & _T_5 | ~_T_5 & _T_3102 : _T_3102;	// sequencer-master.scala:132:52, :184:52
      wire _T_3127 = io_op_bits_active_vfcmp ? _T_2314 & _T_5 | ~_T_5 & _T_3103 : _T_3103;	// sequencer-master.scala:132:52, :184:52
      wire _T_3128 = io_op_bits_active_vfcmp ? _T_2315 & _T_5 | ~_T_5 & _T_3104 : _T_3104;	// sequencer-master.scala:132:52, :184:52
      wire _T_3129 = io_op_bits_active_vfcmp ? _T_2299 & _T_5 | ~_T_5 & _T_3105 : _T_3105;	// sequencer-master.scala:133:52, :185:52
      wire _T_3130 = io_op_bits_active_vfcmp ? _T_2300 & _T_5 | ~_T_5 & _T_3106 : _T_3106;	// sequencer-master.scala:133:52, :185:52
      wire _T_3131 = io_op_bits_active_vfcmp ? _T_2301 & _T_5 | ~_T_5 & _T_3107 : _T_3107;	// sequencer-master.scala:133:52, :185:52
      wire _T_3132 = io_op_bits_active_vfcmp ? _T_2302 & _T_5 | ~_T_5 & _T_3108 : _T_3108;	// sequencer-master.scala:133:52, :185:52
      wire _T_3133 = io_op_bits_active_vfcmp ? _T_2303 & _T_5 | ~_T_5 & _T_3109 : _T_3109;	// sequencer-master.scala:133:52, :185:52
      wire _T_3134 = io_op_bits_active_vfcmp ? _T_2304 & _T_5 | ~_T_5 & _T_3110 : _T_3110;	// sequencer-master.scala:133:52, :185:52
      wire _T_3135 = io_op_bits_active_vfcmp ? _T_2305 & _T_5 | ~_T_5 & _T_3111 : _T_3111;	// sequencer-master.scala:133:52, :185:52
      wire _T_3136 = io_op_bits_active_vfcmp ? _T_2306 & _T_5 | ~_T_5 & _T_3112 : _T_3112;	// sequencer-master.scala:133:52, :185:52
      wire _T_3137 = io_op_bits_active_vfconv ? _T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 & _T_3113 : _T_3113;	// sequencer-master.scala:131:52, :183:52
      wire _T_3138 = io_op_bits_active_vfconv ? _T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 & _T_3114 : _T_3114;	// sequencer-master.scala:131:52, :183:52
      wire _T_3139 = io_op_bits_active_vfconv ? _T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 & _T_3115 : _T_3115;	// sequencer-master.scala:131:52, :183:52
      wire _T_3140 = io_op_bits_active_vfconv ? _T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 & _T_3116 : _T_3116;	// sequencer-master.scala:131:52, :183:52
      wire _T_3141 = io_op_bits_active_vfconv ? _T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 & _T_3117 : _T_3117;	// sequencer-master.scala:131:52, :183:52
      wire _T_3142 = io_op_bits_active_vfconv ? _T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 & _T_3118 : _T_3118;	// sequencer-master.scala:131:52, :183:52
      wire _T_3143 = io_op_bits_active_vfconv ? _T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 & _T_3119 : _T_3119;	// sequencer-master.scala:131:52, :183:52
      wire _T_3144 = io_op_bits_active_vfconv ? _T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 & _T_3120 : _T_3120;	// sequencer-master.scala:131:52, :183:52
      wire _T_3145 = io_op_bits_active_vrpred ? _T_2238 & _T_5 | ~_T_5 & _T_3137 : _T_3137;	// sequencer-master.scala:131:52, :183:52
      wire _T_3146 = io_op_bits_active_vrpred ? _T_2242 & _T_5 | ~_T_5 & _T_3138 : _T_3138;	// sequencer-master.scala:131:52, :183:52
      wire _T_3147 = io_op_bits_active_vrpred ? _T_2246 & _T_5 | ~_T_5 & _T_3139 : _T_3139;	// sequencer-master.scala:131:52, :183:52
      wire _T_3148 = io_op_bits_active_vrpred ? _T_2250 & _T_5 | ~_T_5 & _T_3140 : _T_3140;	// sequencer-master.scala:131:52, :183:52
      wire _T_3149 = io_op_bits_active_vrpred ? _T_2254 & _T_5 | ~_T_5 & _T_3141 : _T_3141;	// sequencer-master.scala:131:52, :183:52
      wire _T_3150 = io_op_bits_active_vrpred ? _T_2258 & _T_5 | ~_T_5 & _T_3142 : _T_3142;	// sequencer-master.scala:131:52, :183:52
      wire _T_3151 = io_op_bits_active_vrpred ? _T_2262 & _T_5 | ~_T_5 & _T_3143 : _T_3143;	// sequencer-master.scala:131:52, :183:52
      wire _T_3152 = io_op_bits_active_vrpred ? _T_2266 & _T_5 | ~_T_5 & _T_3144 : _T_3144;	// sequencer-master.scala:131:52, :183:52
      wire _T_3153 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_5 | ~_T_5 & _T_3121 : _T_3121);	// sequencer-master.scala:132:52, :184:52
      wire _T_3154 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_5 | ~_T_5 & _T_3129 : _T_3129);	// sequencer-master.scala:133:52, :185:52
      wire _T_3155 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_5 | ~_T_5 & _T_3122 : _T_3122);	// sequencer-master.scala:132:52, :184:52
      wire _T_3156 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_5 | ~_T_5 & _T_3130 : _T_3130);	// sequencer-master.scala:133:52, :185:52
      wire _T_3157 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_5 | ~_T_5 & _T_3123 : _T_3123);	// sequencer-master.scala:132:52, :184:52
      wire _T_3158 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_5 | ~_T_5 & _T_3131 : _T_3131);	// sequencer-master.scala:133:52, :185:52
      wire _T_3159 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_5 | ~_T_5 & _T_3124 : _T_3124);	// sequencer-master.scala:132:52, :184:52
      wire _T_3160 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_5 | ~_T_5 & _T_3132 : _T_3132);	// sequencer-master.scala:133:52, :185:52
      wire _T_3161 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_5 | ~_T_5 & _T_3125 : _T_3125);	// sequencer-master.scala:132:52, :184:52
      wire _T_3162 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_5 | ~_T_5 & _T_3133 : _T_3133);	// sequencer-master.scala:133:52, :185:52
      wire _T_3163 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_5 | ~_T_5 & _T_3126 : _T_3126);	// sequencer-master.scala:132:52, :184:52
      wire _T_3164 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_5 | ~_T_5 & _T_3134 : _T_3134);	// sequencer-master.scala:133:52, :185:52
      wire _T_3165 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_5 | ~_T_5 & _T_3127 : _T_3127);	// sequencer-master.scala:132:52, :184:52
      wire _T_3166 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_5 | ~_T_5 & _T_3135 : _T_3135);	// sequencer-master.scala:133:52, :185:52
      wire _T_3167 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_5 | ~_T_5 & _T_3128 : _T_3128);	// sequencer-master.scala:132:52, :184:52
      wire _T_3168 = (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_5 | ~_T_5 & _T_3136 : _T_3136);	// sequencer-master.scala:133:52, :185:52
      wire _T_3169 = io_op_bits_active_vrfirst ? _T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 & _T_3145 : _T_3145;	// sequencer-master.scala:131:52, :183:52
      wire _T_3170 = io_op_bits_active_vrfirst ? _T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 & _T_3146 : _T_3146;	// sequencer-master.scala:131:52, :183:52
      wire _T_3171 = io_op_bits_active_vrfirst ? _T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 & _T_3147 : _T_3147;	// sequencer-master.scala:131:52, :183:52
      wire _T_3172 = io_op_bits_active_vrfirst ? _T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 & _T_3148 : _T_3148;	// sequencer-master.scala:131:52, :183:52
      wire _T_3173 = io_op_bits_active_vrfirst ? _T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 & _T_3149 : _T_3149;	// sequencer-master.scala:131:52, :183:52
      wire _T_3174 = io_op_bits_active_vrfirst ? _T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 & _T_3150 : _T_3150;	// sequencer-master.scala:131:52, :183:52
      wire _T_3175 = io_op_bits_active_vrfirst ? _T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 & _T_3151 : _T_3151;	// sequencer-master.scala:131:52, :183:52
      wire _T_3176 = io_op_bits_active_vrfirst ? _T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 & _T_3152 : _T_3152;	// sequencer-master.scala:131:52, :183:52
      wire _T_3177 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_132 | _T_2279 & _T_292 | _T_2238 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2269 & _T_5 | _T_2238 & _T_5 | ~_T_5 & _T_3169)) : _T_3169;	// sequencer-master.scala:131:52, :183:52
      wire _T_3178 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_133 | _T_2280 & _T_292 | _T_2242 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2270 & _T_5 | _T_2242 & _T_5 | ~_T_5 & _T_3170)) : _T_3170;	// sequencer-master.scala:131:52, :183:52
      wire _T_3179 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_134 | _T_2281 & _T_292 | _T_2246 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2271 & _T_5 | _T_2246 & _T_5 | ~_T_5 & _T_3171)) : _T_3171;	// sequencer-master.scala:131:52, :183:52
      wire _T_3180 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_135 | _T_2282 & _T_292 | _T_2250 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2272 & _T_5 | _T_2250 & _T_5 | ~_T_5 & _T_3172)) : _T_3172;	// sequencer-master.scala:131:52, :183:52
      wire _T_3181 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_136 | _T_2283 & _T_292 | _T_2254 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2273 & _T_5 | _T_2254 & _T_5 | ~_T_5 & _T_3173)) : _T_3173;	// sequencer-master.scala:131:52, :183:52
      wire _T_3182 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_137 | _T_2284 & _T_292 | _T_2258 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2274 & _T_5 | _T_2258 & _T_5 | ~_T_5 & _T_3174)) : _T_3174;	// sequencer-master.scala:131:52, :183:52
      wire _T_3183 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & _T_138 | _T_2285 & _T_292 | _T_2262 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2275 & _T_5 | _T_2262 & _T_5 | ~_T_5 & _T_3175)) : _T_3175;	// sequencer-master.scala:131:52, :183:52
      wire _T_3184 = io_op_bits_active_vamo ? ~_T_315 & (_T_292 & &_T_0 | _T_2286 & _T_292 | _T_2266 & _T_292 |
                ~_T_292 & ~_T_133 & (_T_2276 & _T_5 | _T_2266 & _T_5 | ~_T_5 & _T_3176)) : _T_3176;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3185 = io_op_bits_active_vamo ? _T_2308 & _T_315 | ~_T_315 & ~_T_292 & (_T_2308 & _T_133 | ~_T_133
                & ~_T_5 & _T_3153) : _T_3153;	// sequencer-master.scala:132:52, :184:52
      wire _T_3186 = io_op_bits_active_vamo ? _T_2309 & _T_315 | ~_T_315 & ~_T_292 & (_T_2309 & _T_133 | ~_T_133
                & ~_T_5 & _T_3155) : _T_3155;	// sequencer-master.scala:132:52, :184:52
      wire _T_3187 = io_op_bits_active_vamo ? _T_2310 & _T_315 | ~_T_315 & ~_T_292 & (_T_2310 & _T_133 | ~_T_133
                & ~_T_5 & _T_3157) : _T_3157;	// sequencer-master.scala:132:52, :184:52
      wire _T_3188 = io_op_bits_active_vamo ? _T_2311 & _T_315 | ~_T_315 & ~_T_292 & (_T_2311 & _T_133 | ~_T_133
                & ~_T_5 & _T_3159) : _T_3159;	// sequencer-master.scala:132:52, :184:52
      wire _T_3189 = io_op_bits_active_vamo ? _T_2312 & _T_315 | ~_T_315 & ~_T_292 & (_T_2312 & _T_133 | ~_T_133
                & ~_T_5 & _T_3161) : _T_3161;	// sequencer-master.scala:132:52, :184:52
      wire _T_3190 = io_op_bits_active_vamo ? _T_2313 & _T_315 | ~_T_315 & ~_T_292 & (_T_2313 & _T_133 | ~_T_133
                & ~_T_5 & _T_3163) : _T_3163;	// sequencer-master.scala:132:52, :184:52
      wire _T_3191 = io_op_bits_active_vamo ? _T_2314 & _T_315 | ~_T_315 & ~_T_292 & (_T_2314 & _T_133 | ~_T_133
                & ~_T_5 & _T_3165) : _T_3165;	// sequencer-master.scala:132:52, :184:52
      wire _T_3192 = io_op_bits_active_vamo ? _T_2315 & _T_315 | ~_T_315 & ~_T_292 & (_T_2315 & _T_133 | ~_T_133
                & ~_T_5 & _T_3167) : _T_3167;	// sequencer-master.scala:132:52, :184:52
      wire _T_3193 = io_op_bits_active_vamo ? _T_2299 & _T_315 | ~_T_315 & ~_T_292 & (_T_2299 & _T_133 | ~_T_133
                & ~_T_5 & _T_3154) : _T_3154;	// sequencer-master.scala:133:52, :185:52
      wire _T_3194 = io_op_bits_active_vamo ? _T_2300 & _T_315 | ~_T_315 & ~_T_292 & (_T_2300 & _T_133 | ~_T_133
                & ~_T_5 & _T_3156) : _T_3156;	// sequencer-master.scala:133:52, :185:52
      wire _T_3195 = io_op_bits_active_vamo ? _T_2301 & _T_315 | ~_T_315 & ~_T_292 & (_T_2301 & _T_133 | ~_T_133
                & ~_T_5 & _T_3158) : _T_3158;	// sequencer-master.scala:133:52, :185:52
      wire _T_3196 = io_op_bits_active_vamo ? _T_2302 & _T_315 | ~_T_315 & ~_T_292 & (_T_2302 & _T_133 | ~_T_133
                & ~_T_5 & _T_3160) : _T_3160;	// sequencer-master.scala:133:52, :185:52
      wire _T_3197 = io_op_bits_active_vamo ? _T_2303 & _T_315 | ~_T_315 & ~_T_292 & (_T_2303 & _T_133 | ~_T_133
                & ~_T_5 & _T_3162) : _T_3162;	// sequencer-master.scala:133:52, :185:52
      wire _T_3198 = io_op_bits_active_vamo ? _T_2304 & _T_315 | ~_T_315 & ~_T_292 & (_T_2304 & _T_133 | ~_T_133
                & ~_T_5 & _T_3164) : _T_3164;	// sequencer-master.scala:133:52, :185:52
      wire _T_3199 = io_op_bits_active_vamo ? _T_2305 & _T_315 | ~_T_315 & ~_T_292 & (_T_2305 & _T_133 | ~_T_133
                & ~_T_5 & _T_3166) : _T_3166;	// sequencer-master.scala:133:52, :185:52
      wire _T_3200 = io_op_bits_active_vamo ? _T_2306 & _T_315 | ~_T_315 & ~_T_292 & (_T_2306 & _T_133 | ~_T_133
                & ~_T_5 & _T_3168) : _T_3168;	// sequencer-master.scala:133:52, :185:52
      wire _T_3201 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2279 & _T_5 | _T_2238 & _T_5 | ~_T_5 &
                _T_3177) : _T_3177;	// sequencer-master.scala:131:52, :183:52
      wire _T_3202 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2280 & _T_5 | _T_2242 & _T_5 | ~_T_5 &
                _T_3178) : _T_3178;	// sequencer-master.scala:131:52, :183:52
      wire _T_3203 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2281 & _T_5 | _T_2246 & _T_5 | ~_T_5 &
                _T_3179) : _T_3179;	// sequencer-master.scala:131:52, :183:52
      wire _T_3204 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2282 & _T_5 | _T_2250 & _T_5 | ~_T_5 &
                _T_3180) : _T_3180;	// sequencer-master.scala:131:52, :183:52
      wire _T_3205 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2283 & _T_5 | _T_2254 & _T_5 | ~_T_5 &
                _T_3181) : _T_3181;	// sequencer-master.scala:131:52, :183:52
      wire _T_3206 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2284 & _T_5 | _T_2258 & _T_5 | ~_T_5 &
                _T_3182) : _T_3182;	// sequencer-master.scala:131:52, :183:52
      wire _T_3207 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2285 & _T_5 | _T_2262 & _T_5 | ~_T_5 &
                _T_3183) : _T_3183;	// sequencer-master.scala:131:52, :183:52
      wire _T_3208 = io_op_bits_active_vldx ? ~_T_292 & ~_T_133 & (_T_2286 & _T_5 | _T_2266 & _T_5 | ~_T_5 &
                _T_3184) : _T_3184;	// sequencer-master.scala:131:52, :183:52
      wire _T_3209 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2308 &
                _T_292 | ~_T_292 & (_T_2308 & _T_133 | ~_T_133 & ~_T_5 & _T_3185) : _T_3185);	// sequencer-master.scala:132:52, :184:52
      wire _T_3210 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2299 &
                _T_292 | ~_T_292 & (_T_2299 & _T_133 | ~_T_133 & ~_T_5 & _T_3193) : _T_3193);	// sequencer-master.scala:133:52, :185:52
      wire _T_3211 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2309 &
                _T_292 | ~_T_292 & (_T_2309 & _T_133 | ~_T_133 & ~_T_5 & _T_3186) : _T_3186);	// sequencer-master.scala:132:52, :184:52
      wire _T_3212 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2300 &
                _T_292 | ~_T_292 & (_T_2300 & _T_133 | ~_T_133 & ~_T_5 & _T_3194) : _T_3194);	// sequencer-master.scala:133:52, :185:52
      wire _T_3213 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2310 &
                _T_292 | ~_T_292 & (_T_2310 & _T_133 | ~_T_133 & ~_T_5 & _T_3187) : _T_3187);	// sequencer-master.scala:132:52, :184:52
      wire _T_3214 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2301 &
                _T_292 | ~_T_292 & (_T_2301 & _T_133 | ~_T_133 & ~_T_5 & _T_3195) : _T_3195);	// sequencer-master.scala:133:52, :185:52
      wire _T_3215 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2311 &
                _T_292 | ~_T_292 & (_T_2311 & _T_133 | ~_T_133 & ~_T_5 & _T_3188) : _T_3188);	// sequencer-master.scala:132:52, :184:52
      wire _T_3216 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2302 &
                _T_292 | ~_T_292 & (_T_2302 & _T_133 | ~_T_133 & ~_T_5 & _T_3196) : _T_3196);	// sequencer-master.scala:133:52, :185:52
      wire _T_3217 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2312 &
                _T_292 | ~_T_292 & (_T_2312 & _T_133 | ~_T_133 & ~_T_5 & _T_3189) : _T_3189);	// sequencer-master.scala:132:52, :184:52
      wire _T_3218 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2303 &
                _T_292 | ~_T_292 & (_T_2303 & _T_133 | ~_T_133 & ~_T_5 & _T_3197) : _T_3197);	// sequencer-master.scala:133:52, :185:52
      wire _T_3219 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2313 &
                _T_292 | ~_T_292 & (_T_2313 & _T_133 | ~_T_133 & ~_T_5 & _T_3190) : _T_3190);	// sequencer-master.scala:132:52, :184:52
      wire _T_3220 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2304 &
                _T_292 | ~_T_292 & (_T_2304 & _T_133 | ~_T_133 & ~_T_5 & _T_3198) : _T_3198);	// sequencer-master.scala:133:52, :185:52
      wire _T_3221 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2314 &
                _T_292 | ~_T_292 & (_T_2314 & _T_133 | ~_T_133 & ~_T_5 & _T_3191) : _T_3191);	// sequencer-master.scala:132:52, :184:52
      wire _T_3222 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2305 &
                _T_292 | ~_T_292 & (_T_2305 & _T_133 | ~_T_133 & ~_T_5 & _T_3199) : _T_3199);	// sequencer-master.scala:133:52, :185:52
      wire _T_3223 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2315 &
                _T_292 | ~_T_292 & (_T_2315 & _T_133 | ~_T_133 & ~_T_5 & _T_3192) : _T_3192);	// sequencer-master.scala:132:52, :184:52
      wire _T_3224 = (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vldx ? _T_2306 &
                _T_292 | ~_T_292 & (_T_2306 & _T_133 | ~_T_133 & ~_T_5 & _T_3200) : _T_3200);	// sequencer-master.scala:133:52, :185:52
      wire _T_3225 = io_op_bits_active_vstx ? _T_292 & _T_132 | _T_2299 & _T_292 | _T_2238 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2279 & _T_5 | _T_2238 & _T_5 | ~_T_5 & _T_3201) : _T_3201;	// sequencer-master.scala:131:52, :183:52
      wire _T_3226 = io_op_bits_active_vstx ? _T_292 & _T_133 | _T_2300 & _T_292 | _T_2242 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2280 & _T_5 | _T_2242 & _T_5 | ~_T_5 & _T_3202) : _T_3202;	// sequencer-master.scala:131:52, :183:52
      wire _T_3227 = io_op_bits_active_vstx ? _T_292 & _T_134 | _T_2301 & _T_292 | _T_2246 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2281 & _T_5 | _T_2246 & _T_5 | ~_T_5 & _T_3203) : _T_3203;	// sequencer-master.scala:131:52, :183:52
      wire _T_3228 = io_op_bits_active_vstx ? _T_292 & _T_135 | _T_2302 & _T_292 | _T_2250 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2282 & _T_5 | _T_2250 & _T_5 | ~_T_5 & _T_3204) : _T_3204;	// sequencer-master.scala:131:52, :183:52
      wire _T_3229 = io_op_bits_active_vstx ? _T_292 & _T_136 | _T_2303 & _T_292 | _T_2254 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2283 & _T_5 | _T_2254 & _T_5 | ~_T_5 & _T_3205) : _T_3205;	// sequencer-master.scala:131:52, :183:52
      wire _T_3230 = io_op_bits_active_vstx ? _T_292 & _T_137 | _T_2304 & _T_292 | _T_2258 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2284 & _T_5 | _T_2258 & _T_5 | ~_T_5 & _T_3206) : _T_3206;	// sequencer-master.scala:131:52, :183:52
      wire _T_3231 = io_op_bits_active_vstx ? _T_292 & _T_138 | _T_2305 & _T_292 | _T_2262 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2285 & _T_5 | _T_2262 & _T_5 | ~_T_5 & _T_3207) : _T_3207;	// sequencer-master.scala:131:52, :183:52
      wire _T_3232 = io_op_bits_active_vstx ? _T_292 & &_T_0 | _T_2306 & _T_292 | _T_2266 & _T_292 | ~_T_292 &
                ~_T_133 & (_T_2286 & _T_5 | _T_2266 & _T_5 | ~_T_5 & _T_3208) : _T_3208;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3233 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2238 & _T_5 | ~_T_5 & _T_3225) : _T_3225;	// sequencer-master.scala:131:52, :183:52
      wire _T_3234 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2242 & _T_5 | ~_T_5 & _T_3226) : _T_3226;	// sequencer-master.scala:131:52, :183:52
      wire _T_3235 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2246 & _T_5 | ~_T_5 & _T_3227) : _T_3227;	// sequencer-master.scala:131:52, :183:52
      wire _T_3236 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2250 & _T_5 | ~_T_5 & _T_3228) : _T_3228;	// sequencer-master.scala:131:52, :183:52
      wire _T_3237 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2254 & _T_5 | ~_T_5 & _T_3229) : _T_3229;	// sequencer-master.scala:131:52, :183:52
      wire _T_3238 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2258 & _T_5 | ~_T_5 & _T_3230) : _T_3230;	// sequencer-master.scala:131:52, :183:52
      wire _T_3239 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2262 & _T_5 | ~_T_5 & _T_3231) : _T_3231;	// sequencer-master.scala:131:52, :183:52
      wire _T_3240 = io_op_bits_active_vld ? ~_T_292 & ~_T_133 & (_T_2266 & _T_5 | ~_T_5 & _T_3232) : _T_3232;	// sequencer-master.scala:131:52, :183:52
      wire _T_3241 = io_op_bits_active_vint ? _T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 &
                e_2_raw_0 : e_2_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_3242 = io_op_bits_active_vint ? _T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 &
                e_2_raw_1 : e_2_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_3243 = io_op_bits_active_vint ? _T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 &
                e_2_raw_2 : e_2_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_3244 = io_op_bits_active_vint ? _T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 &
                e_2_raw_3 : e_2_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_3245 = io_op_bits_active_vint ? _T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 &
                e_2_raw_4 : e_2_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_3246 = io_op_bits_active_vint ? _T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 &
                e_2_raw_5 : e_2_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_3247 = io_op_bits_active_vint ? _T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 &
                e_2_raw_6 : e_2_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_3248 = io_op_bits_active_vint ? _T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 &
                e_2_raw_7 : e_2_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_3249 = io_op_bits_active_vint ? _T_2308 & _T_6 | ~_T_6 & e_2_war_0 : e_2_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_3250 = io_op_bits_active_vint ? _T_2309 & _T_6 | ~_T_6 & e_2_war_1 : e_2_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_3251 = io_op_bits_active_vint ? _T_2310 & _T_6 | ~_T_6 & e_2_war_2 : e_2_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_3252 = io_op_bits_active_vint ? _T_2311 & _T_6 | ~_T_6 & e_2_war_3 : e_2_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_3253 = io_op_bits_active_vint ? _T_2312 & _T_6 | ~_T_6 & e_2_war_4 : e_2_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_3254 = io_op_bits_active_vint ? _T_2313 & _T_6 | ~_T_6 & e_2_war_5 : e_2_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_3255 = io_op_bits_active_vint ? _T_2314 & _T_6 | ~_T_6 & e_2_war_6 : e_2_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_3256 = io_op_bits_active_vint ? _T_2315 & _T_6 | ~_T_6 & e_2_war_7 : e_2_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_3257 = io_op_bits_active_vint ? _T_2299 & _T_6 | ~_T_6 & e_2_waw_0 : e_2_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_3258 = io_op_bits_active_vint ? _T_2300 & _T_6 | ~_T_6 & e_2_waw_1 : e_2_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_3259 = io_op_bits_active_vint ? _T_2301 & _T_6 | ~_T_6 & e_2_waw_2 : e_2_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_3260 = io_op_bits_active_vint ? _T_2302 & _T_6 | ~_T_6 & e_2_waw_3 : e_2_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_3261 = io_op_bits_active_vint ? _T_2303 & _T_6 | ~_T_6 & e_2_waw_4 : e_2_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_3262 = io_op_bits_active_vint ? _T_2304 & _T_6 | ~_T_6 & e_2_waw_5 : e_2_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_3263 = io_op_bits_active_vint ? _T_2305 & _T_6 | ~_T_6 & e_2_waw_6 : e_2_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_3264 = io_op_bits_active_vint ? _T_2306 & _T_6 | ~_T_6 & e_2_waw_7 : e_2_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_3265 = io_op_bits_active_vipred ? _T_2289 & _T_6 | _T_2279 & _T_6 | _T_2269 & _T_6 | ~_T_6 &
                _T_3241 : _T_3241;	// sequencer-master.scala:131:52, :183:52
      wire _T_3266 = io_op_bits_active_vipred ? _T_2290 & _T_6 | _T_2280 & _T_6 | _T_2270 & _T_6 | ~_T_6 &
                _T_3242 : _T_3242;	// sequencer-master.scala:131:52, :183:52
      wire _T_3267 = io_op_bits_active_vipred ? _T_2291 & _T_6 | _T_2281 & _T_6 | _T_2271 & _T_6 | ~_T_6 &
                _T_3243 : _T_3243;	// sequencer-master.scala:131:52, :183:52
      wire _T_3268 = io_op_bits_active_vipred ? _T_2292 & _T_6 | _T_2282 & _T_6 | _T_2272 & _T_6 | ~_T_6 &
                _T_3244 : _T_3244;	// sequencer-master.scala:131:52, :183:52
      wire _T_3269 = io_op_bits_active_vipred ? _T_2293 & _T_6 | _T_2283 & _T_6 | _T_2273 & _T_6 | ~_T_6 &
                _T_3245 : _T_3245;	// sequencer-master.scala:131:52, :183:52
      wire _T_3270 = io_op_bits_active_vipred ? _T_2294 & _T_6 | _T_2284 & _T_6 | _T_2274 & _T_6 | ~_T_6 &
                _T_3246 : _T_3246;	// sequencer-master.scala:131:52, :183:52
      wire _T_3271 = io_op_bits_active_vipred ? _T_2295 & _T_6 | _T_2285 & _T_6 | _T_2275 & _T_6 | ~_T_6 &
                _T_3247 : _T_3247;	// sequencer-master.scala:131:52, :183:52
      wire _T_3272 = io_op_bits_active_vipred ? _T_2296 & _T_6 | _T_2286 & _T_6 | _T_2276 & _T_6 | ~_T_6 &
                _T_3248 : _T_3248;	// sequencer-master.scala:131:52, :183:52
      wire _T_3273 = io_op_bits_active_vipred ? _T_2308 & _T_6 | ~_T_6 & _T_3249 : _T_3249;	// sequencer-master.scala:132:52, :184:52
      wire _T_3274 = io_op_bits_active_vipred ? _T_2309 & _T_6 | ~_T_6 & _T_3250 : _T_3250;	// sequencer-master.scala:132:52, :184:52
      wire _T_3275 = io_op_bits_active_vipred ? _T_2310 & _T_6 | ~_T_6 & _T_3251 : _T_3251;	// sequencer-master.scala:132:52, :184:52
      wire _T_3276 = io_op_bits_active_vipred ? _T_2311 & _T_6 | ~_T_6 & _T_3252 : _T_3252;	// sequencer-master.scala:132:52, :184:52
      wire _T_3277 = io_op_bits_active_vipred ? _T_2312 & _T_6 | ~_T_6 & _T_3253 : _T_3253;	// sequencer-master.scala:132:52, :184:52
      wire _T_3278 = io_op_bits_active_vipred ? _T_2313 & _T_6 | ~_T_6 & _T_3254 : _T_3254;	// sequencer-master.scala:132:52, :184:52
      wire _T_3279 = io_op_bits_active_vipred ? _T_2314 & _T_6 | ~_T_6 & _T_3255 : _T_3255;	// sequencer-master.scala:132:52, :184:52
      wire _T_3280 = io_op_bits_active_vipred ? _T_2315 & _T_6 | ~_T_6 & _T_3256 : _T_3256;	// sequencer-master.scala:132:52, :184:52
      wire _T_3281 = io_op_bits_active_vipred ? _T_2299 & _T_6 | ~_T_6 & _T_3257 : _T_3257;	// sequencer-master.scala:133:52, :185:52
      wire _T_3282 = io_op_bits_active_vipred ? _T_2300 & _T_6 | ~_T_6 & _T_3258 : _T_3258;	// sequencer-master.scala:133:52, :185:52
      wire _T_3283 = io_op_bits_active_vipred ? _T_2301 & _T_6 | ~_T_6 & _T_3259 : _T_3259;	// sequencer-master.scala:133:52, :185:52
      wire _T_3284 = io_op_bits_active_vipred ? _T_2302 & _T_6 | ~_T_6 & _T_3260 : _T_3260;	// sequencer-master.scala:133:52, :185:52
      wire _T_3285 = io_op_bits_active_vipred ? _T_2303 & _T_6 | ~_T_6 & _T_3261 : _T_3261;	// sequencer-master.scala:133:52, :185:52
      wire _T_3286 = io_op_bits_active_vipred ? _T_2304 & _T_6 | ~_T_6 & _T_3262 : _T_3262;	// sequencer-master.scala:133:52, :185:52
      wire _T_3287 = io_op_bits_active_vipred ? _T_2305 & _T_6 | ~_T_6 & _T_3263 : _T_3263;	// sequencer-master.scala:133:52, :185:52
      wire _T_3288 = io_op_bits_active_vipred ? _T_2306 & _T_6 | ~_T_6 & _T_3264 : _T_3264;	// sequencer-master.scala:133:52, :185:52
      wire _T_3289 = io_op_bits_active_vimul ? _T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 &
                _T_3265 : _T_3265;	// sequencer-master.scala:131:52, :183:52
      wire _T_3290 = io_op_bits_active_vimul ? _T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 &
                _T_3266 : _T_3266;	// sequencer-master.scala:131:52, :183:52
      wire _T_3291 = io_op_bits_active_vimul ? _T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 &
                _T_3267 : _T_3267;	// sequencer-master.scala:131:52, :183:52
      wire _T_3292 = io_op_bits_active_vimul ? _T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 &
                _T_3268 : _T_3268;	// sequencer-master.scala:131:52, :183:52
      wire _T_3293 = io_op_bits_active_vimul ? _T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 &
                _T_3269 : _T_3269;	// sequencer-master.scala:131:52, :183:52
      wire _T_3294 = io_op_bits_active_vimul ? _T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 &
                _T_3270 : _T_3270;	// sequencer-master.scala:131:52, :183:52
      wire _T_3295 = io_op_bits_active_vimul ? _T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 &
                _T_3271 : _T_3271;	// sequencer-master.scala:131:52, :183:52
      wire _T_3296 = io_op_bits_active_vimul ? _T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 &
                _T_3272 : _T_3272;	// sequencer-master.scala:131:52, :183:52
      wire _T_3297 = io_op_bits_active_vimul ? _T_2308 & _T_6 | ~_T_6 & _T_3273 : _T_3273;	// sequencer-master.scala:132:52, :184:52
      wire _T_3298 = io_op_bits_active_vimul ? _T_2309 & _T_6 | ~_T_6 & _T_3274 : _T_3274;	// sequencer-master.scala:132:52, :184:52
      wire _T_3299 = io_op_bits_active_vimul ? _T_2310 & _T_6 | ~_T_6 & _T_3275 : _T_3275;	// sequencer-master.scala:132:52, :184:52
      wire _T_3300 = io_op_bits_active_vimul ? _T_2311 & _T_6 | ~_T_6 & _T_3276 : _T_3276;	// sequencer-master.scala:132:52, :184:52
      wire _T_3301 = io_op_bits_active_vimul ? _T_2312 & _T_6 | ~_T_6 & _T_3277 : _T_3277;	// sequencer-master.scala:132:52, :184:52
      wire _T_3302 = io_op_bits_active_vimul ? _T_2313 & _T_6 | ~_T_6 & _T_3278 : _T_3278;	// sequencer-master.scala:132:52, :184:52
      wire _T_3303 = io_op_bits_active_vimul ? _T_2314 & _T_6 | ~_T_6 & _T_3279 : _T_3279;	// sequencer-master.scala:132:52, :184:52
      wire _T_3304 = io_op_bits_active_vimul ? _T_2315 & _T_6 | ~_T_6 & _T_3280 : _T_3280;	// sequencer-master.scala:132:52, :184:52
      wire _T_3305 = io_op_bits_active_vimul ? _T_2299 & _T_6 | ~_T_6 & _T_3281 : _T_3281;	// sequencer-master.scala:133:52, :185:52
      wire _T_3306 = io_op_bits_active_vimul ? _T_2300 & _T_6 | ~_T_6 & _T_3282 : _T_3282;	// sequencer-master.scala:133:52, :185:52
      wire _T_3307 = io_op_bits_active_vimul ? _T_2301 & _T_6 | ~_T_6 & _T_3283 : _T_3283;	// sequencer-master.scala:133:52, :185:52
      wire _T_3308 = io_op_bits_active_vimul ? _T_2302 & _T_6 | ~_T_6 & _T_3284 : _T_3284;	// sequencer-master.scala:133:52, :185:52
      wire _T_3309 = io_op_bits_active_vimul ? _T_2303 & _T_6 | ~_T_6 & _T_3285 : _T_3285;	// sequencer-master.scala:133:52, :185:52
      wire _T_3310 = io_op_bits_active_vimul ? _T_2304 & _T_6 | ~_T_6 & _T_3286 : _T_3286;	// sequencer-master.scala:133:52, :185:52
      wire _T_3311 = io_op_bits_active_vimul ? _T_2305 & _T_6 | ~_T_6 & _T_3287 : _T_3287;	// sequencer-master.scala:133:52, :185:52
      wire _T_3312 = io_op_bits_active_vimul ? _T_2306 & _T_6 | ~_T_6 & _T_3288 : _T_3288;	// sequencer-master.scala:133:52, :185:52
      wire _T_3313 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6 |
                ~_T_6 & _T_3289) : _T_3289;	// sequencer-master.scala:131:52, :183:52
      wire _T_3314 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6 |
                ~_T_6 & _T_3290) : _T_3290;	// sequencer-master.scala:131:52, :183:52
      wire _T_3315 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6 |
                ~_T_6 & _T_3291) : _T_3291;	// sequencer-master.scala:131:52, :183:52
      wire _T_3316 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6 |
                ~_T_6 & _T_3292) : _T_3292;	// sequencer-master.scala:131:52, :183:52
      wire _T_3317 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6 |
                ~_T_6 & _T_3293) : _T_3293;	// sequencer-master.scala:131:52, :183:52
      wire _T_3318 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6 |
                ~_T_6 & _T_3294) : _T_3294;	// sequencer-master.scala:131:52, :183:52
      wire _T_3319 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6 |
                ~_T_6 & _T_3295) : _T_3295;	// sequencer-master.scala:131:52, :183:52
      wire _T_3320 = io_op_bits_active_vidiv ? ~_T_134 & (_T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6 |
                ~_T_6 & _T_3296) : _T_3296;	// sequencer-master.scala:131:52, :183:52
      wire _T_3321 = io_op_bits_active_vidiv ? _T_2308 & _T_134 | ~_T_134 & (_T_2308 & _T_6 | ~_T_6 & _T_3297) :
                _T_3297;	// sequencer-master.scala:132:52, :184:52
      wire _T_3322 = io_op_bits_active_vidiv ? _T_2309 & _T_134 | ~_T_134 & (_T_2309 & _T_6 | ~_T_6 & _T_3298) :
                _T_3298;	// sequencer-master.scala:132:52, :184:52
      wire _T_3323 = io_op_bits_active_vidiv ? _T_2310 & _T_134 | ~_T_134 & (_T_2310 & _T_6 | ~_T_6 & _T_3299) :
                _T_3299;	// sequencer-master.scala:132:52, :184:52
      wire _T_3324 = io_op_bits_active_vidiv ? _T_2311 & _T_134 | ~_T_134 & (_T_2311 & _T_6 | ~_T_6 & _T_3300) :
                _T_3300;	// sequencer-master.scala:132:52, :184:52
      wire _T_3325 = io_op_bits_active_vidiv ? _T_2312 & _T_134 | ~_T_134 & (_T_2312 & _T_6 | ~_T_6 & _T_3301) :
                _T_3301;	// sequencer-master.scala:132:52, :184:52
      wire _T_3326 = io_op_bits_active_vidiv ? _T_2313 & _T_134 | ~_T_134 & (_T_2313 & _T_6 | ~_T_6 & _T_3302) :
                _T_3302;	// sequencer-master.scala:132:52, :184:52
      wire _T_3327 = io_op_bits_active_vidiv ? _T_2314 & _T_134 | ~_T_134 & (_T_2314 & _T_6 | ~_T_6 & _T_3303) :
                _T_3303;	// sequencer-master.scala:132:52, :184:52
      wire _T_3328 = io_op_bits_active_vidiv ? _T_2315 & _T_134 | ~_T_134 & (_T_2315 & _T_6 | ~_T_6 & _T_3304) :
                _T_3304;	// sequencer-master.scala:132:52, :184:52
      wire _T_3329 = io_op_bits_active_vidiv ? _T_2299 & _T_134 | ~_T_134 & (_T_2299 & _T_6 | ~_T_6 & _T_3305) :
                _T_3305;	// sequencer-master.scala:133:52, :185:52
      wire _T_3330 = io_op_bits_active_vidiv ? _T_2300 & _T_134 | ~_T_134 & (_T_2300 & _T_6 | ~_T_6 & _T_3306) :
                _T_3306;	// sequencer-master.scala:133:52, :185:52
      wire _T_3331 = io_op_bits_active_vidiv ? _T_2301 & _T_134 | ~_T_134 & (_T_2301 & _T_6 | ~_T_6 & _T_3307) :
                _T_3307;	// sequencer-master.scala:133:52, :185:52
      wire _T_3332 = io_op_bits_active_vidiv ? _T_2302 & _T_134 | ~_T_134 & (_T_2302 & _T_6 | ~_T_6 & _T_3308) :
                _T_3308;	// sequencer-master.scala:133:52, :185:52
      wire _T_3333 = io_op_bits_active_vidiv ? _T_2303 & _T_134 | ~_T_134 & (_T_2303 & _T_6 | ~_T_6 & _T_3309) :
                _T_3309;	// sequencer-master.scala:133:52, :185:52
      wire _T_3334 = io_op_bits_active_vidiv ? _T_2304 & _T_134 | ~_T_134 & (_T_2304 & _T_6 | ~_T_6 & _T_3310) :
                _T_3310;	// sequencer-master.scala:133:52, :185:52
      wire _T_3335 = io_op_bits_active_vidiv ? _T_2305 & _T_134 | ~_T_134 & (_T_2305 & _T_6 | ~_T_6 & _T_3311) :
                _T_3311;	// sequencer-master.scala:133:52, :185:52
      wire _T_3336 = io_op_bits_active_vidiv ? _T_2306 & _T_134 | ~_T_134 & (_T_2306 & _T_6 | ~_T_6 & _T_3312) :
                _T_3312;	// sequencer-master.scala:133:52, :185:52
      wire _T_3337 = io_op_bits_active_vfma ? _T_2289 & _T_6 | _T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6
                | ~_T_6 & _T_3313 : _T_3313;	// sequencer-master.scala:131:52, :183:52
      wire _T_3338 = io_op_bits_active_vfma ? _T_2290 & _T_6 | _T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6
                | ~_T_6 & _T_3314 : _T_3314;	// sequencer-master.scala:131:52, :183:52
      wire _T_3339 = io_op_bits_active_vfma ? _T_2291 & _T_6 | _T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6
                | ~_T_6 & _T_3315 : _T_3315;	// sequencer-master.scala:131:52, :183:52
      wire _T_3340 = io_op_bits_active_vfma ? _T_2292 & _T_6 | _T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6
                | ~_T_6 & _T_3316 : _T_3316;	// sequencer-master.scala:131:52, :183:52
      wire _T_3341 = io_op_bits_active_vfma ? _T_2293 & _T_6 | _T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6
                | ~_T_6 & _T_3317 : _T_3317;	// sequencer-master.scala:131:52, :183:52
      wire _T_3342 = io_op_bits_active_vfma ? _T_2294 & _T_6 | _T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6
                | ~_T_6 & _T_3318 : _T_3318;	// sequencer-master.scala:131:52, :183:52
      wire _T_3343 = io_op_bits_active_vfma ? _T_2295 & _T_6 | _T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6
                | ~_T_6 & _T_3319 : _T_3319;	// sequencer-master.scala:131:52, :183:52
      wire _T_3344 = io_op_bits_active_vfma ? _T_2296 & _T_6 | _T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6
                | ~_T_6 & _T_3320 : _T_3320;	// sequencer-master.scala:131:52, :183:52
      wire _T_3345 = io_op_bits_active_vfma ? _T_2308 & _T_6 | ~_T_6 & _T_3321 : _T_3321;	// sequencer-master.scala:132:52, :184:52
      wire _T_3346 = io_op_bits_active_vfma ? _T_2309 & _T_6 | ~_T_6 & _T_3322 : _T_3322;	// sequencer-master.scala:132:52, :184:52
      wire _T_3347 = io_op_bits_active_vfma ? _T_2310 & _T_6 | ~_T_6 & _T_3323 : _T_3323;	// sequencer-master.scala:132:52, :184:52
      wire _T_3348 = io_op_bits_active_vfma ? _T_2311 & _T_6 | ~_T_6 & _T_3324 : _T_3324;	// sequencer-master.scala:132:52, :184:52
      wire _T_3349 = io_op_bits_active_vfma ? _T_2312 & _T_6 | ~_T_6 & _T_3325 : _T_3325;	// sequencer-master.scala:132:52, :184:52
      wire _T_3350 = io_op_bits_active_vfma ? _T_2313 & _T_6 | ~_T_6 & _T_3326 : _T_3326;	// sequencer-master.scala:132:52, :184:52
      wire _T_3351 = io_op_bits_active_vfma ? _T_2314 & _T_6 | ~_T_6 & _T_3327 : _T_3327;	// sequencer-master.scala:132:52, :184:52
      wire _T_3352 = io_op_bits_active_vfma ? _T_2315 & _T_6 | ~_T_6 & _T_3328 : _T_3328;	// sequencer-master.scala:132:52, :184:52
      wire _T_3353 = io_op_bits_active_vfma ? _T_2299 & _T_6 | ~_T_6 & _T_3329 : _T_3329;	// sequencer-master.scala:133:52, :185:52
      wire _T_3354 = io_op_bits_active_vfma ? _T_2300 & _T_6 | ~_T_6 & _T_3330 : _T_3330;	// sequencer-master.scala:133:52, :185:52
      wire _T_3355 = io_op_bits_active_vfma ? _T_2301 & _T_6 | ~_T_6 & _T_3331 : _T_3331;	// sequencer-master.scala:133:52, :185:52
      wire _T_3356 = io_op_bits_active_vfma ? _T_2302 & _T_6 | ~_T_6 & _T_3332 : _T_3332;	// sequencer-master.scala:133:52, :185:52
      wire _T_3357 = io_op_bits_active_vfma ? _T_2303 & _T_6 | ~_T_6 & _T_3333 : _T_3333;	// sequencer-master.scala:133:52, :185:52
      wire _T_3358 = io_op_bits_active_vfma ? _T_2304 & _T_6 | ~_T_6 & _T_3334 : _T_3334;	// sequencer-master.scala:133:52, :185:52
      wire _T_3359 = io_op_bits_active_vfma ? _T_2305 & _T_6 | ~_T_6 & _T_3335 : _T_3335;	// sequencer-master.scala:133:52, :185:52
      wire _T_3360 = io_op_bits_active_vfma ? _T_2306 & _T_6 | ~_T_6 & _T_3336 : _T_3336;	// sequencer-master.scala:133:52, :185:52
      wire _T_3361 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6 |
                ~_T_6 & _T_3337) : _T_3337;	// sequencer-master.scala:131:52, :183:52
      wire _T_3362 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6 |
                ~_T_6 & _T_3338) : _T_3338;	// sequencer-master.scala:131:52, :183:52
      wire _T_3363 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6 |
                ~_T_6 & _T_3339) : _T_3339;	// sequencer-master.scala:131:52, :183:52
      wire _T_3364 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6 |
                ~_T_6 & _T_3340) : _T_3340;	// sequencer-master.scala:131:52, :183:52
      wire _T_3365 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6 |
                ~_T_6 & _T_3341) : _T_3341;	// sequencer-master.scala:131:52, :183:52
      wire _T_3366 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6 |
                ~_T_6 & _T_3342) : _T_3342;	// sequencer-master.scala:131:52, :183:52
      wire _T_3367 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6 |
                ~_T_6 & _T_3343) : _T_3343;	// sequencer-master.scala:131:52, :183:52
      wire _T_3368 = io_op_bits_active_vfdiv ? ~_T_134 & (_T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6 |
                ~_T_6 & _T_3344) : _T_3344;	// sequencer-master.scala:131:52, :183:52
      wire _T_3369 = io_op_bits_active_vfdiv ? _T_2308 & _T_134 | ~_T_134 & (_T_2308 & _T_6 | ~_T_6 & _T_3345) :
                _T_3345;	// sequencer-master.scala:132:52, :184:52
      wire _T_3370 = io_op_bits_active_vfdiv ? _T_2309 & _T_134 | ~_T_134 & (_T_2309 & _T_6 | ~_T_6 & _T_3346) :
                _T_3346;	// sequencer-master.scala:132:52, :184:52
      wire _T_3371 = io_op_bits_active_vfdiv ? _T_2310 & _T_134 | ~_T_134 & (_T_2310 & _T_6 | ~_T_6 & _T_3347) :
                _T_3347;	// sequencer-master.scala:132:52, :184:52
      wire _T_3372 = io_op_bits_active_vfdiv ? _T_2311 & _T_134 | ~_T_134 & (_T_2311 & _T_6 | ~_T_6 & _T_3348) :
                _T_3348;	// sequencer-master.scala:132:52, :184:52
      wire _T_3373 = io_op_bits_active_vfdiv ? _T_2312 & _T_134 | ~_T_134 & (_T_2312 & _T_6 | ~_T_6 & _T_3349) :
                _T_3349;	// sequencer-master.scala:132:52, :184:52
      wire _T_3374 = io_op_bits_active_vfdiv ? _T_2313 & _T_134 | ~_T_134 & (_T_2313 & _T_6 | ~_T_6 & _T_3350) :
                _T_3350;	// sequencer-master.scala:132:52, :184:52
      wire _T_3375 = io_op_bits_active_vfdiv ? _T_2314 & _T_134 | ~_T_134 & (_T_2314 & _T_6 | ~_T_6 & _T_3351) :
                _T_3351;	// sequencer-master.scala:132:52, :184:52
      wire _T_3376 = io_op_bits_active_vfdiv ? _T_2315 & _T_134 | ~_T_134 & (_T_2315 & _T_6 | ~_T_6 & _T_3352) :
                _T_3352;	// sequencer-master.scala:132:52, :184:52
      wire _T_3377 = io_op_bits_active_vfdiv ? _T_2299 & _T_134 | ~_T_134 & (_T_2299 & _T_6 | ~_T_6 & _T_3353) :
                _T_3353;	// sequencer-master.scala:133:52, :185:52
      wire _T_3378 = io_op_bits_active_vfdiv ? _T_2300 & _T_134 | ~_T_134 & (_T_2300 & _T_6 | ~_T_6 & _T_3354) :
                _T_3354;	// sequencer-master.scala:133:52, :185:52
      wire _T_3379 = io_op_bits_active_vfdiv ? _T_2301 & _T_134 | ~_T_134 & (_T_2301 & _T_6 | ~_T_6 & _T_3355) :
                _T_3355;	// sequencer-master.scala:133:52, :185:52
      wire _T_3380 = io_op_bits_active_vfdiv ? _T_2302 & _T_134 | ~_T_134 & (_T_2302 & _T_6 | ~_T_6 & _T_3356) :
                _T_3356;	// sequencer-master.scala:133:52, :185:52
      wire _T_3381 = io_op_bits_active_vfdiv ? _T_2303 & _T_134 | ~_T_134 & (_T_2303 & _T_6 | ~_T_6 & _T_3357) :
                _T_3357;	// sequencer-master.scala:133:52, :185:52
      wire _T_3382 = io_op_bits_active_vfdiv ? _T_2304 & _T_134 | ~_T_134 & (_T_2304 & _T_6 | ~_T_6 & _T_3358) :
                _T_3358;	// sequencer-master.scala:133:52, :185:52
      wire _T_3383 = io_op_bits_active_vfdiv ? _T_2305 & _T_134 | ~_T_134 & (_T_2305 & _T_6 | ~_T_6 & _T_3359) :
                _T_3359;	// sequencer-master.scala:133:52, :185:52
      wire _T_3384 = io_op_bits_active_vfdiv ? _T_2306 & _T_134 | ~_T_134 & (_T_2306 & _T_6 | ~_T_6 & _T_3360) :
                _T_3360;	// sequencer-master.scala:133:52, :185:52
      wire _T_3385 = io_op_bits_active_vfcmp ? _T_2279 & _T_6 | _T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 &
                _T_3361 : _T_3361;	// sequencer-master.scala:131:52, :183:52
      wire _T_3386 = io_op_bits_active_vfcmp ? _T_2280 & _T_6 | _T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 &
                _T_3362 : _T_3362;	// sequencer-master.scala:131:52, :183:52
      wire _T_3387 = io_op_bits_active_vfcmp ? _T_2281 & _T_6 | _T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 &
                _T_3363 : _T_3363;	// sequencer-master.scala:131:52, :183:52
      wire _T_3388 = io_op_bits_active_vfcmp ? _T_2282 & _T_6 | _T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 &
                _T_3364 : _T_3364;	// sequencer-master.scala:131:52, :183:52
      wire _T_3389 = io_op_bits_active_vfcmp ? _T_2283 & _T_6 | _T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 &
                _T_3365 : _T_3365;	// sequencer-master.scala:131:52, :183:52
      wire _T_3390 = io_op_bits_active_vfcmp ? _T_2284 & _T_6 | _T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 &
                _T_3366 : _T_3366;	// sequencer-master.scala:131:52, :183:52
      wire _T_3391 = io_op_bits_active_vfcmp ? _T_2285 & _T_6 | _T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 &
                _T_3367 : _T_3367;	// sequencer-master.scala:131:52, :183:52
      wire _T_3392 = io_op_bits_active_vfcmp ? _T_2286 & _T_6 | _T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 &
                _T_3368 : _T_3368;	// sequencer-master.scala:131:52, :183:52
      wire _T_3393 = io_op_bits_active_vfcmp ? _T_2308 & _T_6 | ~_T_6 & _T_3369 : _T_3369;	// sequencer-master.scala:132:52, :184:52
      wire _T_3394 = io_op_bits_active_vfcmp ? _T_2309 & _T_6 | ~_T_6 & _T_3370 : _T_3370;	// sequencer-master.scala:132:52, :184:52
      wire _T_3395 = io_op_bits_active_vfcmp ? _T_2310 & _T_6 | ~_T_6 & _T_3371 : _T_3371;	// sequencer-master.scala:132:52, :184:52
      wire _T_3396 = io_op_bits_active_vfcmp ? _T_2311 & _T_6 | ~_T_6 & _T_3372 : _T_3372;	// sequencer-master.scala:132:52, :184:52
      wire _T_3397 = io_op_bits_active_vfcmp ? _T_2312 & _T_6 | ~_T_6 & _T_3373 : _T_3373;	// sequencer-master.scala:132:52, :184:52
      wire _T_3398 = io_op_bits_active_vfcmp ? _T_2313 & _T_6 | ~_T_6 & _T_3374 : _T_3374;	// sequencer-master.scala:132:52, :184:52
      wire _T_3399 = io_op_bits_active_vfcmp ? _T_2314 & _T_6 | ~_T_6 & _T_3375 : _T_3375;	// sequencer-master.scala:132:52, :184:52
      wire _T_3400 = io_op_bits_active_vfcmp ? _T_2315 & _T_6 | ~_T_6 & _T_3376 : _T_3376;	// sequencer-master.scala:132:52, :184:52
      wire _T_3401 = io_op_bits_active_vfcmp ? _T_2299 & _T_6 | ~_T_6 & _T_3377 : _T_3377;	// sequencer-master.scala:133:52, :185:52
      wire _T_3402 = io_op_bits_active_vfcmp ? _T_2300 & _T_6 | ~_T_6 & _T_3378 : _T_3378;	// sequencer-master.scala:133:52, :185:52
      wire _T_3403 = io_op_bits_active_vfcmp ? _T_2301 & _T_6 | ~_T_6 & _T_3379 : _T_3379;	// sequencer-master.scala:133:52, :185:52
      wire _T_3404 = io_op_bits_active_vfcmp ? _T_2302 & _T_6 | ~_T_6 & _T_3380 : _T_3380;	// sequencer-master.scala:133:52, :185:52
      wire _T_3405 = io_op_bits_active_vfcmp ? _T_2303 & _T_6 | ~_T_6 & _T_3381 : _T_3381;	// sequencer-master.scala:133:52, :185:52
      wire _T_3406 = io_op_bits_active_vfcmp ? _T_2304 & _T_6 | ~_T_6 & _T_3382 : _T_3382;	// sequencer-master.scala:133:52, :185:52
      wire _T_3407 = io_op_bits_active_vfcmp ? _T_2305 & _T_6 | ~_T_6 & _T_3383 : _T_3383;	// sequencer-master.scala:133:52, :185:52
      wire _T_3408 = io_op_bits_active_vfcmp ? _T_2306 & _T_6 | ~_T_6 & _T_3384 : _T_3384;	// sequencer-master.scala:133:52, :185:52
      wire _T_3409 = io_op_bits_active_vfconv ? _T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 & _T_3385 : _T_3385;	// sequencer-master.scala:131:52, :183:52
      wire _T_3410 = io_op_bits_active_vfconv ? _T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 & _T_3386 : _T_3386;	// sequencer-master.scala:131:52, :183:52
      wire _T_3411 = io_op_bits_active_vfconv ? _T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 & _T_3387 : _T_3387;	// sequencer-master.scala:131:52, :183:52
      wire _T_3412 = io_op_bits_active_vfconv ? _T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 & _T_3388 : _T_3388;	// sequencer-master.scala:131:52, :183:52
      wire _T_3413 = io_op_bits_active_vfconv ? _T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 & _T_3389 : _T_3389;	// sequencer-master.scala:131:52, :183:52
      wire _T_3414 = io_op_bits_active_vfconv ? _T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 & _T_3390 : _T_3390;	// sequencer-master.scala:131:52, :183:52
      wire _T_3415 = io_op_bits_active_vfconv ? _T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 & _T_3391 : _T_3391;	// sequencer-master.scala:131:52, :183:52
      wire _T_3416 = io_op_bits_active_vfconv ? _T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 & _T_3392 : _T_3392;	// sequencer-master.scala:131:52, :183:52
      wire _T_3417 = io_op_bits_active_vrpred ? _T_2238 & _T_6 | ~_T_6 & _T_3409 : _T_3409;	// sequencer-master.scala:131:52, :183:52
      wire _T_3418 = io_op_bits_active_vrpred ? _T_2242 & _T_6 | ~_T_6 & _T_3410 : _T_3410;	// sequencer-master.scala:131:52, :183:52
      wire _T_3419 = io_op_bits_active_vrpred ? _T_2246 & _T_6 | ~_T_6 & _T_3411 : _T_3411;	// sequencer-master.scala:131:52, :183:52
      wire _T_3420 = io_op_bits_active_vrpred ? _T_2250 & _T_6 | ~_T_6 & _T_3412 : _T_3412;	// sequencer-master.scala:131:52, :183:52
      wire _T_3421 = io_op_bits_active_vrpred ? _T_2254 & _T_6 | ~_T_6 & _T_3413 : _T_3413;	// sequencer-master.scala:131:52, :183:52
      wire _T_3422 = io_op_bits_active_vrpred ? _T_2258 & _T_6 | ~_T_6 & _T_3414 : _T_3414;	// sequencer-master.scala:131:52, :183:52
      wire _T_3423 = io_op_bits_active_vrpred ? _T_2262 & _T_6 | ~_T_6 & _T_3415 : _T_3415;	// sequencer-master.scala:131:52, :183:52
      wire _T_3424 = io_op_bits_active_vrpred ? _T_2266 & _T_6 | ~_T_6 & _T_3416 : _T_3416;	// sequencer-master.scala:131:52, :183:52
      wire _T_3425 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_6 | ~_T_6 & _T_3393 : _T_3393);	// sequencer-master.scala:132:52, :184:52
      wire _T_3426 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_6 | ~_T_6 & _T_3401 : _T_3401);	// sequencer-master.scala:133:52, :185:52
      wire _T_3427 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_6 | ~_T_6 & _T_3394 : _T_3394);	// sequencer-master.scala:132:52, :184:52
      wire _T_3428 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_6 | ~_T_6 & _T_3402 : _T_3402);	// sequencer-master.scala:133:52, :185:52
      wire _T_3429 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_6 | ~_T_6 & _T_3395 : _T_3395);	// sequencer-master.scala:132:52, :184:52
      wire _T_3430 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_6 | ~_T_6 & _T_3403 : _T_3403);	// sequencer-master.scala:133:52, :185:52
      wire _T_3431 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_6 | ~_T_6 & _T_3396 : _T_3396);	// sequencer-master.scala:132:52, :184:52
      wire _T_3432 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_6 | ~_T_6 & _T_3404 : _T_3404);	// sequencer-master.scala:133:52, :185:52
      wire _T_3433 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_6 | ~_T_6 & _T_3397 : _T_3397);	// sequencer-master.scala:132:52, :184:52
      wire _T_3434 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_6 | ~_T_6 & _T_3405 : _T_3405);	// sequencer-master.scala:133:52, :185:52
      wire _T_3435 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_6 | ~_T_6 & _T_3398 : _T_3398);	// sequencer-master.scala:132:52, :184:52
      wire _T_3436 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_6 | ~_T_6 & _T_3406 : _T_3406);	// sequencer-master.scala:133:52, :185:52
      wire _T_3437 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_6 | ~_T_6 & _T_3399 : _T_3399);	// sequencer-master.scala:132:52, :184:52
      wire _T_3438 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_6 | ~_T_6 & _T_3407 : _T_3407);	// sequencer-master.scala:133:52, :185:52
      wire _T_3439 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_6 | ~_T_6 & _T_3400 : _T_3400);	// sequencer-master.scala:132:52, :184:52
      wire _T_3440 = (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_6 | ~_T_6 & _T_3408 : _T_3408);	// sequencer-master.scala:133:52, :185:52
      wire _T_3441 = io_op_bits_active_vrfirst ? _T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 & _T_3417 : _T_3417;	// sequencer-master.scala:131:52, :183:52
      wire _T_3442 = io_op_bits_active_vrfirst ? _T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 & _T_3418 : _T_3418;	// sequencer-master.scala:131:52, :183:52
      wire _T_3443 = io_op_bits_active_vrfirst ? _T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 & _T_3419 : _T_3419;	// sequencer-master.scala:131:52, :183:52
      wire _T_3444 = io_op_bits_active_vrfirst ? _T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 & _T_3420 : _T_3420;	// sequencer-master.scala:131:52, :183:52
      wire _T_3445 = io_op_bits_active_vrfirst ? _T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 & _T_3421 : _T_3421;	// sequencer-master.scala:131:52, :183:52
      wire _T_3446 = io_op_bits_active_vrfirst ? _T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 & _T_3422 : _T_3422;	// sequencer-master.scala:131:52, :183:52
      wire _T_3447 = io_op_bits_active_vrfirst ? _T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 & _T_3423 : _T_3423;	// sequencer-master.scala:131:52, :183:52
      wire _T_3448 = io_op_bits_active_vrfirst ? _T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 & _T_3424 : _T_3424;	// sequencer-master.scala:131:52, :183:52
      wire _T_3449 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_132 | _T_2279 & _T_293 | _T_2238 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2269 & _T_6 | _T_2238 & _T_6 | ~_T_6 & _T_3441)) : _T_3441;	// sequencer-master.scala:131:52, :183:52
      wire _T_3450 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_133 | _T_2280 & _T_293 | _T_2242 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2270 & _T_6 | _T_2242 & _T_6 | ~_T_6 & _T_3442)) : _T_3442;	// sequencer-master.scala:131:52, :183:52
      wire _T_3451 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_134 | _T_2281 & _T_293 | _T_2246 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2271 & _T_6 | _T_2246 & _T_6 | ~_T_6 & _T_3443)) : _T_3443;	// sequencer-master.scala:131:52, :183:52
      wire _T_3452 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_135 | _T_2282 & _T_293 | _T_2250 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2272 & _T_6 | _T_2250 & _T_6 | ~_T_6 & _T_3444)) : _T_3444;	// sequencer-master.scala:131:52, :183:52
      wire _T_3453 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_136 | _T_2283 & _T_293 | _T_2254 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2273 & _T_6 | _T_2254 & _T_6 | ~_T_6 & _T_3445)) : _T_3445;	// sequencer-master.scala:131:52, :183:52
      wire _T_3454 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_137 | _T_2284 & _T_293 | _T_2258 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2274 & _T_6 | _T_2258 & _T_6 | ~_T_6 & _T_3446)) : _T_3446;	// sequencer-master.scala:131:52, :183:52
      wire _T_3455 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & _T_138 | _T_2285 & _T_293 | _T_2262 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2275 & _T_6 | _T_2262 & _T_6 | ~_T_6 & _T_3447)) : _T_3447;	// sequencer-master.scala:131:52, :183:52
      wire _T_3456 = io_op_bits_active_vamo ? ~_T_316 & (_T_293 & &_T_0 | _T_2286 & _T_293 | _T_2266 & _T_293 |
                ~_T_293 & ~_T_134 & (_T_2276 & _T_6 | _T_2266 & _T_6 | ~_T_6 & _T_3448)) : _T_3448;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3457 = io_op_bits_active_vamo ? _T_2308 & _T_316 | ~_T_316 & ~_T_293 & (_T_2308 & _T_134 | ~_T_134
                & ~_T_6 & _T_3425) : _T_3425;	// sequencer-master.scala:132:52, :184:52
      wire _T_3458 = io_op_bits_active_vamo ? _T_2309 & _T_316 | ~_T_316 & ~_T_293 & (_T_2309 & _T_134 | ~_T_134
                & ~_T_6 & _T_3427) : _T_3427;	// sequencer-master.scala:132:52, :184:52
      wire _T_3459 = io_op_bits_active_vamo ? _T_2310 & _T_316 | ~_T_316 & ~_T_293 & (_T_2310 & _T_134 | ~_T_134
                & ~_T_6 & _T_3429) : _T_3429;	// sequencer-master.scala:132:52, :184:52
      wire _T_3460 = io_op_bits_active_vamo ? _T_2311 & _T_316 | ~_T_316 & ~_T_293 & (_T_2311 & _T_134 | ~_T_134
                & ~_T_6 & _T_3431) : _T_3431;	// sequencer-master.scala:132:52, :184:52
      wire _T_3461 = io_op_bits_active_vamo ? _T_2312 & _T_316 | ~_T_316 & ~_T_293 & (_T_2312 & _T_134 | ~_T_134
                & ~_T_6 & _T_3433) : _T_3433;	// sequencer-master.scala:132:52, :184:52
      wire _T_3462 = io_op_bits_active_vamo ? _T_2313 & _T_316 | ~_T_316 & ~_T_293 & (_T_2313 & _T_134 | ~_T_134
                & ~_T_6 & _T_3435) : _T_3435;	// sequencer-master.scala:132:52, :184:52
      wire _T_3463 = io_op_bits_active_vamo ? _T_2314 & _T_316 | ~_T_316 & ~_T_293 & (_T_2314 & _T_134 | ~_T_134
                & ~_T_6 & _T_3437) : _T_3437;	// sequencer-master.scala:132:52, :184:52
      wire _T_3464 = io_op_bits_active_vamo ? _T_2315 & _T_316 | ~_T_316 & ~_T_293 & (_T_2315 & _T_134 | ~_T_134
                & ~_T_6 & _T_3439) : _T_3439;	// sequencer-master.scala:132:52, :184:52
      wire _T_3465 = io_op_bits_active_vamo ? _T_2299 & _T_316 | ~_T_316 & ~_T_293 & (_T_2299 & _T_134 | ~_T_134
                & ~_T_6 & _T_3426) : _T_3426;	// sequencer-master.scala:133:52, :185:52
      wire _T_3466 = io_op_bits_active_vamo ? _T_2300 & _T_316 | ~_T_316 & ~_T_293 & (_T_2300 & _T_134 | ~_T_134
                & ~_T_6 & _T_3428) : _T_3428;	// sequencer-master.scala:133:52, :185:52
      wire _T_3467 = io_op_bits_active_vamo ? _T_2301 & _T_316 | ~_T_316 & ~_T_293 & (_T_2301 & _T_134 | ~_T_134
                & ~_T_6 & _T_3430) : _T_3430;	// sequencer-master.scala:133:52, :185:52
      wire _T_3468 = io_op_bits_active_vamo ? _T_2302 & _T_316 | ~_T_316 & ~_T_293 & (_T_2302 & _T_134 | ~_T_134
                & ~_T_6 & _T_3432) : _T_3432;	// sequencer-master.scala:133:52, :185:52
      wire _T_3469 = io_op_bits_active_vamo ? _T_2303 & _T_316 | ~_T_316 & ~_T_293 & (_T_2303 & _T_134 | ~_T_134
                & ~_T_6 & _T_3434) : _T_3434;	// sequencer-master.scala:133:52, :185:52
      wire _T_3470 = io_op_bits_active_vamo ? _T_2304 & _T_316 | ~_T_316 & ~_T_293 & (_T_2304 & _T_134 | ~_T_134
                & ~_T_6 & _T_3436) : _T_3436;	// sequencer-master.scala:133:52, :185:52
      wire _T_3471 = io_op_bits_active_vamo ? _T_2305 & _T_316 | ~_T_316 & ~_T_293 & (_T_2305 & _T_134 | ~_T_134
                & ~_T_6 & _T_3438) : _T_3438;	// sequencer-master.scala:133:52, :185:52
      wire _T_3472 = io_op_bits_active_vamo ? _T_2306 & _T_316 | ~_T_316 & ~_T_293 & (_T_2306 & _T_134 | ~_T_134
                & ~_T_6 & _T_3440) : _T_3440;	// sequencer-master.scala:133:52, :185:52
      wire _T_3473 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2279 & _T_6 | _T_2238 & _T_6 | ~_T_6 &
                _T_3449) : _T_3449;	// sequencer-master.scala:131:52, :183:52
      wire _T_3474 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2280 & _T_6 | _T_2242 & _T_6 | ~_T_6 &
                _T_3450) : _T_3450;	// sequencer-master.scala:131:52, :183:52
      wire _T_3475 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2281 & _T_6 | _T_2246 & _T_6 | ~_T_6 &
                _T_3451) : _T_3451;	// sequencer-master.scala:131:52, :183:52
      wire _T_3476 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2282 & _T_6 | _T_2250 & _T_6 | ~_T_6 &
                _T_3452) : _T_3452;	// sequencer-master.scala:131:52, :183:52
      wire _T_3477 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2283 & _T_6 | _T_2254 & _T_6 | ~_T_6 &
                _T_3453) : _T_3453;	// sequencer-master.scala:131:52, :183:52
      wire _T_3478 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2284 & _T_6 | _T_2258 & _T_6 | ~_T_6 &
                _T_3454) : _T_3454;	// sequencer-master.scala:131:52, :183:52
      wire _T_3479 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2285 & _T_6 | _T_2262 & _T_6 | ~_T_6 &
                _T_3455) : _T_3455;	// sequencer-master.scala:131:52, :183:52
      wire _T_3480 = io_op_bits_active_vldx ? ~_T_293 & ~_T_134 & (_T_2286 & _T_6 | _T_2266 & _T_6 | ~_T_6 &
                _T_3456) : _T_3456;	// sequencer-master.scala:131:52, :183:52
      wire _T_3481 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2308 &
                _T_293 | ~_T_293 & (_T_2308 & _T_134 | ~_T_134 & ~_T_6 & _T_3457) : _T_3457);	// sequencer-master.scala:132:52, :184:52
      wire _T_3482 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2299 &
                _T_293 | ~_T_293 & (_T_2299 & _T_134 | ~_T_134 & ~_T_6 & _T_3465) : _T_3465);	// sequencer-master.scala:133:52, :185:52
      wire _T_3483 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2309 &
                _T_293 | ~_T_293 & (_T_2309 & _T_134 | ~_T_134 & ~_T_6 & _T_3458) : _T_3458);	// sequencer-master.scala:132:52, :184:52
      wire _T_3484 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2300 &
                _T_293 | ~_T_293 & (_T_2300 & _T_134 | ~_T_134 & ~_T_6 & _T_3466) : _T_3466);	// sequencer-master.scala:133:52, :185:52
      wire _T_3485 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2310 &
                _T_293 | ~_T_293 & (_T_2310 & _T_134 | ~_T_134 & ~_T_6 & _T_3459) : _T_3459);	// sequencer-master.scala:132:52, :184:52
      wire _T_3486 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2301 &
                _T_293 | ~_T_293 & (_T_2301 & _T_134 | ~_T_134 & ~_T_6 & _T_3467) : _T_3467);	// sequencer-master.scala:133:52, :185:52
      wire _T_3487 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2311 &
                _T_293 | ~_T_293 & (_T_2311 & _T_134 | ~_T_134 & ~_T_6 & _T_3460) : _T_3460);	// sequencer-master.scala:132:52, :184:52
      wire _T_3488 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2302 &
                _T_293 | ~_T_293 & (_T_2302 & _T_134 | ~_T_134 & ~_T_6 & _T_3468) : _T_3468);	// sequencer-master.scala:133:52, :185:52
      wire _T_3489 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2312 &
                _T_293 | ~_T_293 & (_T_2312 & _T_134 | ~_T_134 & ~_T_6 & _T_3461) : _T_3461);	// sequencer-master.scala:132:52, :184:52
      wire _T_3490 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2303 &
                _T_293 | ~_T_293 & (_T_2303 & _T_134 | ~_T_134 & ~_T_6 & _T_3469) : _T_3469);	// sequencer-master.scala:133:52, :185:52
      wire _T_3491 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2313 &
                _T_293 | ~_T_293 & (_T_2313 & _T_134 | ~_T_134 & ~_T_6 & _T_3462) : _T_3462);	// sequencer-master.scala:132:52, :184:52
      wire _T_3492 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2304 &
                _T_293 | ~_T_293 & (_T_2304 & _T_134 | ~_T_134 & ~_T_6 & _T_3470) : _T_3470);	// sequencer-master.scala:133:52, :185:52
      wire _T_3493 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2314 &
                _T_293 | ~_T_293 & (_T_2314 & _T_134 | ~_T_134 & ~_T_6 & _T_3463) : _T_3463);	// sequencer-master.scala:132:52, :184:52
      wire _T_3494 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2305 &
                _T_293 | ~_T_293 & (_T_2305 & _T_134 | ~_T_134 & ~_T_6 & _T_3471) : _T_3471);	// sequencer-master.scala:133:52, :185:52
      wire _T_3495 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2315 &
                _T_293 | ~_T_293 & (_T_2315 & _T_134 | ~_T_134 & ~_T_6 & _T_3464) : _T_3464);	// sequencer-master.scala:132:52, :184:52
      wire _T_3496 = (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vldx ? _T_2306 &
                _T_293 | ~_T_293 & (_T_2306 & _T_134 | ~_T_134 & ~_T_6 & _T_3472) : _T_3472);	// sequencer-master.scala:133:52, :185:52
      wire _T_3497 = io_op_bits_active_vstx ? _T_293 & _T_132 | _T_2299 & _T_293 | _T_2238 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2279 & _T_6 | _T_2238 & _T_6 | ~_T_6 & _T_3473) : _T_3473;	// sequencer-master.scala:131:52, :183:52
      wire _T_3498 = io_op_bits_active_vstx ? _T_293 & _T_133 | _T_2300 & _T_293 | _T_2242 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2280 & _T_6 | _T_2242 & _T_6 | ~_T_6 & _T_3474) : _T_3474;	// sequencer-master.scala:131:52, :183:52
      wire _T_3499 = io_op_bits_active_vstx ? _T_293 & _T_134 | _T_2301 & _T_293 | _T_2246 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2281 & _T_6 | _T_2246 & _T_6 | ~_T_6 & _T_3475) : _T_3475;	// sequencer-master.scala:131:52, :183:52
      wire _T_3500 = io_op_bits_active_vstx ? _T_293 & _T_135 | _T_2302 & _T_293 | _T_2250 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2282 & _T_6 | _T_2250 & _T_6 | ~_T_6 & _T_3476) : _T_3476;	// sequencer-master.scala:131:52, :183:52
      wire _T_3501 = io_op_bits_active_vstx ? _T_293 & _T_136 | _T_2303 & _T_293 | _T_2254 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2283 & _T_6 | _T_2254 & _T_6 | ~_T_6 & _T_3477) : _T_3477;	// sequencer-master.scala:131:52, :183:52
      wire _T_3502 = io_op_bits_active_vstx ? _T_293 & _T_137 | _T_2304 & _T_293 | _T_2258 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2284 & _T_6 | _T_2258 & _T_6 | ~_T_6 & _T_3478) : _T_3478;	// sequencer-master.scala:131:52, :183:52
      wire _T_3503 = io_op_bits_active_vstx ? _T_293 & _T_138 | _T_2305 & _T_293 | _T_2262 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2285 & _T_6 | _T_2262 & _T_6 | ~_T_6 & _T_3479) : _T_3479;	// sequencer-master.scala:131:52, :183:52
      wire _T_3504 = io_op_bits_active_vstx ? _T_293 & &_T_0 | _T_2306 & _T_293 | _T_2266 & _T_293 | ~_T_293 &
                ~_T_134 & (_T_2286 & _T_6 | _T_2266 & _T_6 | ~_T_6 & _T_3480) : _T_3480;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3505 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2238 & _T_6 | ~_T_6 & _T_3497) : _T_3497;	// sequencer-master.scala:131:52, :183:52
      wire _T_3506 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2242 & _T_6 | ~_T_6 & _T_3498) : _T_3498;	// sequencer-master.scala:131:52, :183:52
      wire _T_3507 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2246 & _T_6 | ~_T_6 & _T_3499) : _T_3499;	// sequencer-master.scala:131:52, :183:52
      wire _T_3508 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2250 & _T_6 | ~_T_6 & _T_3500) : _T_3500;	// sequencer-master.scala:131:52, :183:52
      wire _T_3509 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2254 & _T_6 | ~_T_6 & _T_3501) : _T_3501;	// sequencer-master.scala:131:52, :183:52
      wire _T_3510 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2258 & _T_6 | ~_T_6 & _T_3502) : _T_3502;	// sequencer-master.scala:131:52, :183:52
      wire _T_3511 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2262 & _T_6 | ~_T_6 & _T_3503) : _T_3503;	// sequencer-master.scala:131:52, :183:52
      wire _T_3512 = io_op_bits_active_vld ? ~_T_293 & ~_T_134 & (_T_2266 & _T_6 | ~_T_6 & _T_3504) : _T_3504;	// sequencer-master.scala:131:52, :183:52
      wire _T_3513 = io_op_bits_active_vint ? _T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 &
                e_3_raw_0 : e_3_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_3514 = io_op_bits_active_vint ? _T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 &
                e_3_raw_1 : e_3_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_3515 = io_op_bits_active_vint ? _T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 &
                e_3_raw_2 : e_3_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_3516 = io_op_bits_active_vint ? _T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 &
                e_3_raw_3 : e_3_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_3517 = io_op_bits_active_vint ? _T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 &
                e_3_raw_4 : e_3_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_3518 = io_op_bits_active_vint ? _T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 &
                e_3_raw_5 : e_3_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_3519 = io_op_bits_active_vint ? _T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 &
                e_3_raw_6 : e_3_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_3520 = io_op_bits_active_vint ? _T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 &
                e_3_raw_7 : e_3_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_3521 = io_op_bits_active_vint ? _T_2308 & _T_7 | ~_T_7 & e_3_war_0 : e_3_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_3522 = io_op_bits_active_vint ? _T_2309 & _T_7 | ~_T_7 & e_3_war_1 : e_3_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_3523 = io_op_bits_active_vint ? _T_2310 & _T_7 | ~_T_7 & e_3_war_2 : e_3_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_3524 = io_op_bits_active_vint ? _T_2311 & _T_7 | ~_T_7 & e_3_war_3 : e_3_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_3525 = io_op_bits_active_vint ? _T_2312 & _T_7 | ~_T_7 & e_3_war_4 : e_3_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_3526 = io_op_bits_active_vint ? _T_2313 & _T_7 | ~_T_7 & e_3_war_5 : e_3_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_3527 = io_op_bits_active_vint ? _T_2314 & _T_7 | ~_T_7 & e_3_war_6 : e_3_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_3528 = io_op_bits_active_vint ? _T_2315 & _T_7 | ~_T_7 & e_3_war_7 : e_3_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_3529 = io_op_bits_active_vint ? _T_2299 & _T_7 | ~_T_7 & e_3_waw_0 : e_3_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_3530 = io_op_bits_active_vint ? _T_2300 & _T_7 | ~_T_7 & e_3_waw_1 : e_3_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_3531 = io_op_bits_active_vint ? _T_2301 & _T_7 | ~_T_7 & e_3_waw_2 : e_3_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_3532 = io_op_bits_active_vint ? _T_2302 & _T_7 | ~_T_7 & e_3_waw_3 : e_3_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_3533 = io_op_bits_active_vint ? _T_2303 & _T_7 | ~_T_7 & e_3_waw_4 : e_3_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_3534 = io_op_bits_active_vint ? _T_2304 & _T_7 | ~_T_7 & e_3_waw_5 : e_3_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_3535 = io_op_bits_active_vint ? _T_2305 & _T_7 | ~_T_7 & e_3_waw_6 : e_3_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_3536 = io_op_bits_active_vint ? _T_2306 & _T_7 | ~_T_7 & e_3_waw_7 : e_3_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_3537 = io_op_bits_active_vipred ? _T_2289 & _T_7 | _T_2279 & _T_7 | _T_2269 & _T_7 | ~_T_7 &
                _T_3513 : _T_3513;	// sequencer-master.scala:131:52, :183:52
      wire _T_3538 = io_op_bits_active_vipred ? _T_2290 & _T_7 | _T_2280 & _T_7 | _T_2270 & _T_7 | ~_T_7 &
                _T_3514 : _T_3514;	// sequencer-master.scala:131:52, :183:52
      wire _T_3539 = io_op_bits_active_vipred ? _T_2291 & _T_7 | _T_2281 & _T_7 | _T_2271 & _T_7 | ~_T_7 &
                _T_3515 : _T_3515;	// sequencer-master.scala:131:52, :183:52
      wire _T_3540 = io_op_bits_active_vipred ? _T_2292 & _T_7 | _T_2282 & _T_7 | _T_2272 & _T_7 | ~_T_7 &
                _T_3516 : _T_3516;	// sequencer-master.scala:131:52, :183:52
      wire _T_3541 = io_op_bits_active_vipred ? _T_2293 & _T_7 | _T_2283 & _T_7 | _T_2273 & _T_7 | ~_T_7 &
                _T_3517 : _T_3517;	// sequencer-master.scala:131:52, :183:52
      wire _T_3542 = io_op_bits_active_vipred ? _T_2294 & _T_7 | _T_2284 & _T_7 | _T_2274 & _T_7 | ~_T_7 &
                _T_3518 : _T_3518;	// sequencer-master.scala:131:52, :183:52
      wire _T_3543 = io_op_bits_active_vipred ? _T_2295 & _T_7 | _T_2285 & _T_7 | _T_2275 & _T_7 | ~_T_7 &
                _T_3519 : _T_3519;	// sequencer-master.scala:131:52, :183:52
      wire _T_3544 = io_op_bits_active_vipred ? _T_2296 & _T_7 | _T_2286 & _T_7 | _T_2276 & _T_7 | ~_T_7 &
                _T_3520 : _T_3520;	// sequencer-master.scala:131:52, :183:52
      wire _T_3545 = io_op_bits_active_vipred ? _T_2308 & _T_7 | ~_T_7 & _T_3521 : _T_3521;	// sequencer-master.scala:132:52, :184:52
      wire _T_3546 = io_op_bits_active_vipred ? _T_2309 & _T_7 | ~_T_7 & _T_3522 : _T_3522;	// sequencer-master.scala:132:52, :184:52
      wire _T_3547 = io_op_bits_active_vipred ? _T_2310 & _T_7 | ~_T_7 & _T_3523 : _T_3523;	// sequencer-master.scala:132:52, :184:52
      wire _T_3548 = io_op_bits_active_vipred ? _T_2311 & _T_7 | ~_T_7 & _T_3524 : _T_3524;	// sequencer-master.scala:132:52, :184:52
      wire _T_3549 = io_op_bits_active_vipred ? _T_2312 & _T_7 | ~_T_7 & _T_3525 : _T_3525;	// sequencer-master.scala:132:52, :184:52
      wire _T_3550 = io_op_bits_active_vipred ? _T_2313 & _T_7 | ~_T_7 & _T_3526 : _T_3526;	// sequencer-master.scala:132:52, :184:52
      wire _T_3551 = io_op_bits_active_vipred ? _T_2314 & _T_7 | ~_T_7 & _T_3527 : _T_3527;	// sequencer-master.scala:132:52, :184:52
      wire _T_3552 = io_op_bits_active_vipred ? _T_2315 & _T_7 | ~_T_7 & _T_3528 : _T_3528;	// sequencer-master.scala:132:52, :184:52
      wire _T_3553 = io_op_bits_active_vipred ? _T_2299 & _T_7 | ~_T_7 & _T_3529 : _T_3529;	// sequencer-master.scala:133:52, :185:52
      wire _T_3554 = io_op_bits_active_vipred ? _T_2300 & _T_7 | ~_T_7 & _T_3530 : _T_3530;	// sequencer-master.scala:133:52, :185:52
      wire _T_3555 = io_op_bits_active_vipred ? _T_2301 & _T_7 | ~_T_7 & _T_3531 : _T_3531;	// sequencer-master.scala:133:52, :185:52
      wire _T_3556 = io_op_bits_active_vipred ? _T_2302 & _T_7 | ~_T_7 & _T_3532 : _T_3532;	// sequencer-master.scala:133:52, :185:52
      wire _T_3557 = io_op_bits_active_vipred ? _T_2303 & _T_7 | ~_T_7 & _T_3533 : _T_3533;	// sequencer-master.scala:133:52, :185:52
      wire _T_3558 = io_op_bits_active_vipred ? _T_2304 & _T_7 | ~_T_7 & _T_3534 : _T_3534;	// sequencer-master.scala:133:52, :185:52
      wire _T_3559 = io_op_bits_active_vipred ? _T_2305 & _T_7 | ~_T_7 & _T_3535 : _T_3535;	// sequencer-master.scala:133:52, :185:52
      wire _T_3560 = io_op_bits_active_vipred ? _T_2306 & _T_7 | ~_T_7 & _T_3536 : _T_3536;	// sequencer-master.scala:133:52, :185:52
      wire _T_3561 = io_op_bits_active_vimul ? _T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 &
                _T_3537 : _T_3537;	// sequencer-master.scala:131:52, :183:52
      wire _T_3562 = io_op_bits_active_vimul ? _T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 &
                _T_3538 : _T_3538;	// sequencer-master.scala:131:52, :183:52
      wire _T_3563 = io_op_bits_active_vimul ? _T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 &
                _T_3539 : _T_3539;	// sequencer-master.scala:131:52, :183:52
      wire _T_3564 = io_op_bits_active_vimul ? _T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 &
                _T_3540 : _T_3540;	// sequencer-master.scala:131:52, :183:52
      wire _T_3565 = io_op_bits_active_vimul ? _T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 &
                _T_3541 : _T_3541;	// sequencer-master.scala:131:52, :183:52
      wire _T_3566 = io_op_bits_active_vimul ? _T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 &
                _T_3542 : _T_3542;	// sequencer-master.scala:131:52, :183:52
      wire _T_3567 = io_op_bits_active_vimul ? _T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 &
                _T_3543 : _T_3543;	// sequencer-master.scala:131:52, :183:52
      wire _T_3568 = io_op_bits_active_vimul ? _T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 &
                _T_3544 : _T_3544;	// sequencer-master.scala:131:52, :183:52
      wire _T_3569 = io_op_bits_active_vimul ? _T_2308 & _T_7 | ~_T_7 & _T_3545 : _T_3545;	// sequencer-master.scala:132:52, :184:52
      wire _T_3570 = io_op_bits_active_vimul ? _T_2309 & _T_7 | ~_T_7 & _T_3546 : _T_3546;	// sequencer-master.scala:132:52, :184:52
      wire _T_3571 = io_op_bits_active_vimul ? _T_2310 & _T_7 | ~_T_7 & _T_3547 : _T_3547;	// sequencer-master.scala:132:52, :184:52
      wire _T_3572 = io_op_bits_active_vimul ? _T_2311 & _T_7 | ~_T_7 & _T_3548 : _T_3548;	// sequencer-master.scala:132:52, :184:52
      wire _T_3573 = io_op_bits_active_vimul ? _T_2312 & _T_7 | ~_T_7 & _T_3549 : _T_3549;	// sequencer-master.scala:132:52, :184:52
      wire _T_3574 = io_op_bits_active_vimul ? _T_2313 & _T_7 | ~_T_7 & _T_3550 : _T_3550;	// sequencer-master.scala:132:52, :184:52
      wire _T_3575 = io_op_bits_active_vimul ? _T_2314 & _T_7 | ~_T_7 & _T_3551 : _T_3551;	// sequencer-master.scala:132:52, :184:52
      wire _T_3576 = io_op_bits_active_vimul ? _T_2315 & _T_7 | ~_T_7 & _T_3552 : _T_3552;	// sequencer-master.scala:132:52, :184:52
      wire _T_3577 = io_op_bits_active_vimul ? _T_2299 & _T_7 | ~_T_7 & _T_3553 : _T_3553;	// sequencer-master.scala:133:52, :185:52
      wire _T_3578 = io_op_bits_active_vimul ? _T_2300 & _T_7 | ~_T_7 & _T_3554 : _T_3554;	// sequencer-master.scala:133:52, :185:52
      wire _T_3579 = io_op_bits_active_vimul ? _T_2301 & _T_7 | ~_T_7 & _T_3555 : _T_3555;	// sequencer-master.scala:133:52, :185:52
      wire _T_3580 = io_op_bits_active_vimul ? _T_2302 & _T_7 | ~_T_7 & _T_3556 : _T_3556;	// sequencer-master.scala:133:52, :185:52
      wire _T_3581 = io_op_bits_active_vimul ? _T_2303 & _T_7 | ~_T_7 & _T_3557 : _T_3557;	// sequencer-master.scala:133:52, :185:52
      wire _T_3582 = io_op_bits_active_vimul ? _T_2304 & _T_7 | ~_T_7 & _T_3558 : _T_3558;	// sequencer-master.scala:133:52, :185:52
      wire _T_3583 = io_op_bits_active_vimul ? _T_2305 & _T_7 | ~_T_7 & _T_3559 : _T_3559;	// sequencer-master.scala:133:52, :185:52
      wire _T_3584 = io_op_bits_active_vimul ? _T_2306 & _T_7 | ~_T_7 & _T_3560 : _T_3560;	// sequencer-master.scala:133:52, :185:52
      wire _T_3585 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7 |
                ~_T_7 & _T_3561) : _T_3561;	// sequencer-master.scala:131:52, :183:52
      wire _T_3586 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7 |
                ~_T_7 & _T_3562) : _T_3562;	// sequencer-master.scala:131:52, :183:52
      wire _T_3587 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7 |
                ~_T_7 & _T_3563) : _T_3563;	// sequencer-master.scala:131:52, :183:52
      wire _T_3588 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7 |
                ~_T_7 & _T_3564) : _T_3564;	// sequencer-master.scala:131:52, :183:52
      wire _T_3589 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7 |
                ~_T_7 & _T_3565) : _T_3565;	// sequencer-master.scala:131:52, :183:52
      wire _T_3590 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7 |
                ~_T_7 & _T_3566) : _T_3566;	// sequencer-master.scala:131:52, :183:52
      wire _T_3591 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7 |
                ~_T_7 & _T_3567) : _T_3567;	// sequencer-master.scala:131:52, :183:52
      wire _T_3592 = io_op_bits_active_vidiv ? ~_T_135 & (_T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7 |
                ~_T_7 & _T_3568) : _T_3568;	// sequencer-master.scala:131:52, :183:52
      wire _T_3593 = io_op_bits_active_vidiv ? _T_2308 & _T_135 | ~_T_135 & (_T_2308 & _T_7 | ~_T_7 & _T_3569) :
                _T_3569;	// sequencer-master.scala:132:52, :184:52
      wire _T_3594 = io_op_bits_active_vidiv ? _T_2309 & _T_135 | ~_T_135 & (_T_2309 & _T_7 | ~_T_7 & _T_3570) :
                _T_3570;	// sequencer-master.scala:132:52, :184:52
      wire _T_3595 = io_op_bits_active_vidiv ? _T_2310 & _T_135 | ~_T_135 & (_T_2310 & _T_7 | ~_T_7 & _T_3571) :
                _T_3571;	// sequencer-master.scala:132:52, :184:52
      wire _T_3596 = io_op_bits_active_vidiv ? _T_2311 & _T_135 | ~_T_135 & (_T_2311 & _T_7 | ~_T_7 & _T_3572) :
                _T_3572;	// sequencer-master.scala:132:52, :184:52
      wire _T_3597 = io_op_bits_active_vidiv ? _T_2312 & _T_135 | ~_T_135 & (_T_2312 & _T_7 | ~_T_7 & _T_3573) :
                _T_3573;	// sequencer-master.scala:132:52, :184:52
      wire _T_3598 = io_op_bits_active_vidiv ? _T_2313 & _T_135 | ~_T_135 & (_T_2313 & _T_7 | ~_T_7 & _T_3574) :
                _T_3574;	// sequencer-master.scala:132:52, :184:52
      wire _T_3599 = io_op_bits_active_vidiv ? _T_2314 & _T_135 | ~_T_135 & (_T_2314 & _T_7 | ~_T_7 & _T_3575) :
                _T_3575;	// sequencer-master.scala:132:52, :184:52
      wire _T_3600 = io_op_bits_active_vidiv ? _T_2315 & _T_135 | ~_T_135 & (_T_2315 & _T_7 | ~_T_7 & _T_3576) :
                _T_3576;	// sequencer-master.scala:132:52, :184:52
      wire _T_3601 = io_op_bits_active_vidiv ? _T_2299 & _T_135 | ~_T_135 & (_T_2299 & _T_7 | ~_T_7 & _T_3577) :
                _T_3577;	// sequencer-master.scala:133:52, :185:52
      wire _T_3602 = io_op_bits_active_vidiv ? _T_2300 & _T_135 | ~_T_135 & (_T_2300 & _T_7 | ~_T_7 & _T_3578) :
                _T_3578;	// sequencer-master.scala:133:52, :185:52
      wire _T_3603 = io_op_bits_active_vidiv ? _T_2301 & _T_135 | ~_T_135 & (_T_2301 & _T_7 | ~_T_7 & _T_3579) :
                _T_3579;	// sequencer-master.scala:133:52, :185:52
      wire _T_3604 = io_op_bits_active_vidiv ? _T_2302 & _T_135 | ~_T_135 & (_T_2302 & _T_7 | ~_T_7 & _T_3580) :
                _T_3580;	// sequencer-master.scala:133:52, :185:52
      wire _T_3605 = io_op_bits_active_vidiv ? _T_2303 & _T_135 | ~_T_135 & (_T_2303 & _T_7 | ~_T_7 & _T_3581) :
                _T_3581;	// sequencer-master.scala:133:52, :185:52
      wire _T_3606 = io_op_bits_active_vidiv ? _T_2304 & _T_135 | ~_T_135 & (_T_2304 & _T_7 | ~_T_7 & _T_3582) :
                _T_3582;	// sequencer-master.scala:133:52, :185:52
      wire _T_3607 = io_op_bits_active_vidiv ? _T_2305 & _T_135 | ~_T_135 & (_T_2305 & _T_7 | ~_T_7 & _T_3583) :
                _T_3583;	// sequencer-master.scala:133:52, :185:52
      wire _T_3608 = io_op_bits_active_vidiv ? _T_2306 & _T_135 | ~_T_135 & (_T_2306 & _T_7 | ~_T_7 & _T_3584) :
                _T_3584;	// sequencer-master.scala:133:52, :185:52
      wire _T_3609 = io_op_bits_active_vfma ? _T_2289 & _T_7 | _T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7
                | ~_T_7 & _T_3585 : _T_3585;	// sequencer-master.scala:131:52, :183:52
      wire _T_3610 = io_op_bits_active_vfma ? _T_2290 & _T_7 | _T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7
                | ~_T_7 & _T_3586 : _T_3586;	// sequencer-master.scala:131:52, :183:52
      wire _T_3611 = io_op_bits_active_vfma ? _T_2291 & _T_7 | _T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7
                | ~_T_7 & _T_3587 : _T_3587;	// sequencer-master.scala:131:52, :183:52
      wire _T_3612 = io_op_bits_active_vfma ? _T_2292 & _T_7 | _T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7
                | ~_T_7 & _T_3588 : _T_3588;	// sequencer-master.scala:131:52, :183:52
      wire _T_3613 = io_op_bits_active_vfma ? _T_2293 & _T_7 | _T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7
                | ~_T_7 & _T_3589 : _T_3589;	// sequencer-master.scala:131:52, :183:52
      wire _T_3614 = io_op_bits_active_vfma ? _T_2294 & _T_7 | _T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7
                | ~_T_7 & _T_3590 : _T_3590;	// sequencer-master.scala:131:52, :183:52
      wire _T_3615 = io_op_bits_active_vfma ? _T_2295 & _T_7 | _T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7
                | ~_T_7 & _T_3591 : _T_3591;	// sequencer-master.scala:131:52, :183:52
      wire _T_3616 = io_op_bits_active_vfma ? _T_2296 & _T_7 | _T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7
                | ~_T_7 & _T_3592 : _T_3592;	// sequencer-master.scala:131:52, :183:52
      wire _T_3617 = io_op_bits_active_vfma ? _T_2308 & _T_7 | ~_T_7 & _T_3593 : _T_3593;	// sequencer-master.scala:132:52, :184:52
      wire _T_3618 = io_op_bits_active_vfma ? _T_2309 & _T_7 | ~_T_7 & _T_3594 : _T_3594;	// sequencer-master.scala:132:52, :184:52
      wire _T_3619 = io_op_bits_active_vfma ? _T_2310 & _T_7 | ~_T_7 & _T_3595 : _T_3595;	// sequencer-master.scala:132:52, :184:52
      wire _T_3620 = io_op_bits_active_vfma ? _T_2311 & _T_7 | ~_T_7 & _T_3596 : _T_3596;	// sequencer-master.scala:132:52, :184:52
      wire _T_3621 = io_op_bits_active_vfma ? _T_2312 & _T_7 | ~_T_7 & _T_3597 : _T_3597;	// sequencer-master.scala:132:52, :184:52
      wire _T_3622 = io_op_bits_active_vfma ? _T_2313 & _T_7 | ~_T_7 & _T_3598 : _T_3598;	// sequencer-master.scala:132:52, :184:52
      wire _T_3623 = io_op_bits_active_vfma ? _T_2314 & _T_7 | ~_T_7 & _T_3599 : _T_3599;	// sequencer-master.scala:132:52, :184:52
      wire _T_3624 = io_op_bits_active_vfma ? _T_2315 & _T_7 | ~_T_7 & _T_3600 : _T_3600;	// sequencer-master.scala:132:52, :184:52
      wire _T_3625 = io_op_bits_active_vfma ? _T_2299 & _T_7 | ~_T_7 & _T_3601 : _T_3601;	// sequencer-master.scala:133:52, :185:52
      wire _T_3626 = io_op_bits_active_vfma ? _T_2300 & _T_7 | ~_T_7 & _T_3602 : _T_3602;	// sequencer-master.scala:133:52, :185:52
      wire _T_3627 = io_op_bits_active_vfma ? _T_2301 & _T_7 | ~_T_7 & _T_3603 : _T_3603;	// sequencer-master.scala:133:52, :185:52
      wire _T_3628 = io_op_bits_active_vfma ? _T_2302 & _T_7 | ~_T_7 & _T_3604 : _T_3604;	// sequencer-master.scala:133:52, :185:52
      wire _T_3629 = io_op_bits_active_vfma ? _T_2303 & _T_7 | ~_T_7 & _T_3605 : _T_3605;	// sequencer-master.scala:133:52, :185:52
      wire _T_3630 = io_op_bits_active_vfma ? _T_2304 & _T_7 | ~_T_7 & _T_3606 : _T_3606;	// sequencer-master.scala:133:52, :185:52
      wire _T_3631 = io_op_bits_active_vfma ? _T_2305 & _T_7 | ~_T_7 & _T_3607 : _T_3607;	// sequencer-master.scala:133:52, :185:52
      wire _T_3632 = io_op_bits_active_vfma ? _T_2306 & _T_7 | ~_T_7 & _T_3608 : _T_3608;	// sequencer-master.scala:133:52, :185:52
      wire _T_3633 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7 |
                ~_T_7 & _T_3609) : _T_3609;	// sequencer-master.scala:131:52, :183:52
      wire _T_3634 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7 |
                ~_T_7 & _T_3610) : _T_3610;	// sequencer-master.scala:131:52, :183:52
      wire _T_3635 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7 |
                ~_T_7 & _T_3611) : _T_3611;	// sequencer-master.scala:131:52, :183:52
      wire _T_3636 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7 |
                ~_T_7 & _T_3612) : _T_3612;	// sequencer-master.scala:131:52, :183:52
      wire _T_3637 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7 |
                ~_T_7 & _T_3613) : _T_3613;	// sequencer-master.scala:131:52, :183:52
      wire _T_3638 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7 |
                ~_T_7 & _T_3614) : _T_3614;	// sequencer-master.scala:131:52, :183:52
      wire _T_3639 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7 |
                ~_T_7 & _T_3615) : _T_3615;	// sequencer-master.scala:131:52, :183:52
      wire _T_3640 = io_op_bits_active_vfdiv ? ~_T_135 & (_T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7 |
                ~_T_7 & _T_3616) : _T_3616;	// sequencer-master.scala:131:52, :183:52
      wire _T_3641 = io_op_bits_active_vfdiv ? _T_2308 & _T_135 | ~_T_135 & (_T_2308 & _T_7 | ~_T_7 & _T_3617) :
                _T_3617;	// sequencer-master.scala:132:52, :184:52
      wire _T_3642 = io_op_bits_active_vfdiv ? _T_2309 & _T_135 | ~_T_135 & (_T_2309 & _T_7 | ~_T_7 & _T_3618) :
                _T_3618;	// sequencer-master.scala:132:52, :184:52
      wire _T_3643 = io_op_bits_active_vfdiv ? _T_2310 & _T_135 | ~_T_135 & (_T_2310 & _T_7 | ~_T_7 & _T_3619) :
                _T_3619;	// sequencer-master.scala:132:52, :184:52
      wire _T_3644 = io_op_bits_active_vfdiv ? _T_2311 & _T_135 | ~_T_135 & (_T_2311 & _T_7 | ~_T_7 & _T_3620) :
                _T_3620;	// sequencer-master.scala:132:52, :184:52
      wire _T_3645 = io_op_bits_active_vfdiv ? _T_2312 & _T_135 | ~_T_135 & (_T_2312 & _T_7 | ~_T_7 & _T_3621) :
                _T_3621;	// sequencer-master.scala:132:52, :184:52
      wire _T_3646 = io_op_bits_active_vfdiv ? _T_2313 & _T_135 | ~_T_135 & (_T_2313 & _T_7 | ~_T_7 & _T_3622) :
                _T_3622;	// sequencer-master.scala:132:52, :184:52
      wire _T_3647 = io_op_bits_active_vfdiv ? _T_2314 & _T_135 | ~_T_135 & (_T_2314 & _T_7 | ~_T_7 & _T_3623) :
                _T_3623;	// sequencer-master.scala:132:52, :184:52
      wire _T_3648 = io_op_bits_active_vfdiv ? _T_2315 & _T_135 | ~_T_135 & (_T_2315 & _T_7 | ~_T_7 & _T_3624) :
                _T_3624;	// sequencer-master.scala:132:52, :184:52
      wire _T_3649 = io_op_bits_active_vfdiv ? _T_2299 & _T_135 | ~_T_135 & (_T_2299 & _T_7 | ~_T_7 & _T_3625) :
                _T_3625;	// sequencer-master.scala:133:52, :185:52
      wire _T_3650 = io_op_bits_active_vfdiv ? _T_2300 & _T_135 | ~_T_135 & (_T_2300 & _T_7 | ~_T_7 & _T_3626) :
                _T_3626;	// sequencer-master.scala:133:52, :185:52
      wire _T_3651 = io_op_bits_active_vfdiv ? _T_2301 & _T_135 | ~_T_135 & (_T_2301 & _T_7 | ~_T_7 & _T_3627) :
                _T_3627;	// sequencer-master.scala:133:52, :185:52
      wire _T_3652 = io_op_bits_active_vfdiv ? _T_2302 & _T_135 | ~_T_135 & (_T_2302 & _T_7 | ~_T_7 & _T_3628) :
                _T_3628;	// sequencer-master.scala:133:52, :185:52
      wire _T_3653 = io_op_bits_active_vfdiv ? _T_2303 & _T_135 | ~_T_135 & (_T_2303 & _T_7 | ~_T_7 & _T_3629) :
                _T_3629;	// sequencer-master.scala:133:52, :185:52
      wire _T_3654 = io_op_bits_active_vfdiv ? _T_2304 & _T_135 | ~_T_135 & (_T_2304 & _T_7 | ~_T_7 & _T_3630) :
                _T_3630;	// sequencer-master.scala:133:52, :185:52
      wire _T_3655 = io_op_bits_active_vfdiv ? _T_2305 & _T_135 | ~_T_135 & (_T_2305 & _T_7 | ~_T_7 & _T_3631) :
                _T_3631;	// sequencer-master.scala:133:52, :185:52
      wire _T_3656 = io_op_bits_active_vfdiv ? _T_2306 & _T_135 | ~_T_135 & (_T_2306 & _T_7 | ~_T_7 & _T_3632) :
                _T_3632;	// sequencer-master.scala:133:52, :185:52
      wire _T_3657 = io_op_bits_active_vfcmp ? _T_2279 & _T_7 | _T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 &
                _T_3633 : _T_3633;	// sequencer-master.scala:131:52, :183:52
      wire _T_3658 = io_op_bits_active_vfcmp ? _T_2280 & _T_7 | _T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 &
                _T_3634 : _T_3634;	// sequencer-master.scala:131:52, :183:52
      wire _T_3659 = io_op_bits_active_vfcmp ? _T_2281 & _T_7 | _T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 &
                _T_3635 : _T_3635;	// sequencer-master.scala:131:52, :183:52
      wire _T_3660 = io_op_bits_active_vfcmp ? _T_2282 & _T_7 | _T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 &
                _T_3636 : _T_3636;	// sequencer-master.scala:131:52, :183:52
      wire _T_3661 = io_op_bits_active_vfcmp ? _T_2283 & _T_7 | _T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 &
                _T_3637 : _T_3637;	// sequencer-master.scala:131:52, :183:52
      wire _T_3662 = io_op_bits_active_vfcmp ? _T_2284 & _T_7 | _T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 &
                _T_3638 : _T_3638;	// sequencer-master.scala:131:52, :183:52
      wire _T_3663 = io_op_bits_active_vfcmp ? _T_2285 & _T_7 | _T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 &
                _T_3639 : _T_3639;	// sequencer-master.scala:131:52, :183:52
      wire _T_3664 = io_op_bits_active_vfcmp ? _T_2286 & _T_7 | _T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 &
                _T_3640 : _T_3640;	// sequencer-master.scala:131:52, :183:52
      wire _T_3665 = io_op_bits_active_vfcmp ? _T_2308 & _T_7 | ~_T_7 & _T_3641 : _T_3641;	// sequencer-master.scala:132:52, :184:52
      wire _T_3666 = io_op_bits_active_vfcmp ? _T_2309 & _T_7 | ~_T_7 & _T_3642 : _T_3642;	// sequencer-master.scala:132:52, :184:52
      wire _T_3667 = io_op_bits_active_vfcmp ? _T_2310 & _T_7 | ~_T_7 & _T_3643 : _T_3643;	// sequencer-master.scala:132:52, :184:52
      wire _T_3668 = io_op_bits_active_vfcmp ? _T_2311 & _T_7 | ~_T_7 & _T_3644 : _T_3644;	// sequencer-master.scala:132:52, :184:52
      wire _T_3669 = io_op_bits_active_vfcmp ? _T_2312 & _T_7 | ~_T_7 & _T_3645 : _T_3645;	// sequencer-master.scala:132:52, :184:52
      wire _T_3670 = io_op_bits_active_vfcmp ? _T_2313 & _T_7 | ~_T_7 & _T_3646 : _T_3646;	// sequencer-master.scala:132:52, :184:52
      wire _T_3671 = io_op_bits_active_vfcmp ? _T_2314 & _T_7 | ~_T_7 & _T_3647 : _T_3647;	// sequencer-master.scala:132:52, :184:52
      wire _T_3672 = io_op_bits_active_vfcmp ? _T_2315 & _T_7 | ~_T_7 & _T_3648 : _T_3648;	// sequencer-master.scala:132:52, :184:52
      wire _T_3673 = io_op_bits_active_vfcmp ? _T_2299 & _T_7 | ~_T_7 & _T_3649 : _T_3649;	// sequencer-master.scala:133:52, :185:52
      wire _T_3674 = io_op_bits_active_vfcmp ? _T_2300 & _T_7 | ~_T_7 & _T_3650 : _T_3650;	// sequencer-master.scala:133:52, :185:52
      wire _T_3675 = io_op_bits_active_vfcmp ? _T_2301 & _T_7 | ~_T_7 & _T_3651 : _T_3651;	// sequencer-master.scala:133:52, :185:52
      wire _T_3676 = io_op_bits_active_vfcmp ? _T_2302 & _T_7 | ~_T_7 & _T_3652 : _T_3652;	// sequencer-master.scala:133:52, :185:52
      wire _T_3677 = io_op_bits_active_vfcmp ? _T_2303 & _T_7 | ~_T_7 & _T_3653 : _T_3653;	// sequencer-master.scala:133:52, :185:52
      wire _T_3678 = io_op_bits_active_vfcmp ? _T_2304 & _T_7 | ~_T_7 & _T_3654 : _T_3654;	// sequencer-master.scala:133:52, :185:52
      wire _T_3679 = io_op_bits_active_vfcmp ? _T_2305 & _T_7 | ~_T_7 & _T_3655 : _T_3655;	// sequencer-master.scala:133:52, :185:52
      wire _T_3680 = io_op_bits_active_vfcmp ? _T_2306 & _T_7 | ~_T_7 & _T_3656 : _T_3656;	// sequencer-master.scala:133:52, :185:52
      wire _T_3681 = io_op_bits_active_vfconv ? _T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 & _T_3657 : _T_3657;	// sequencer-master.scala:131:52, :183:52
      wire _T_3682 = io_op_bits_active_vfconv ? _T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 & _T_3658 : _T_3658;	// sequencer-master.scala:131:52, :183:52
      wire _T_3683 = io_op_bits_active_vfconv ? _T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 & _T_3659 : _T_3659;	// sequencer-master.scala:131:52, :183:52
      wire _T_3684 = io_op_bits_active_vfconv ? _T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 & _T_3660 : _T_3660;	// sequencer-master.scala:131:52, :183:52
      wire _T_3685 = io_op_bits_active_vfconv ? _T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 & _T_3661 : _T_3661;	// sequencer-master.scala:131:52, :183:52
      wire _T_3686 = io_op_bits_active_vfconv ? _T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 & _T_3662 : _T_3662;	// sequencer-master.scala:131:52, :183:52
      wire _T_3687 = io_op_bits_active_vfconv ? _T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 & _T_3663 : _T_3663;	// sequencer-master.scala:131:52, :183:52
      wire _T_3688 = io_op_bits_active_vfconv ? _T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 & _T_3664 : _T_3664;	// sequencer-master.scala:131:52, :183:52
      wire _T_3689 = io_op_bits_active_vrpred ? _T_2238 & _T_7 | ~_T_7 & _T_3681 : _T_3681;	// sequencer-master.scala:131:52, :183:52
      wire _T_3690 = io_op_bits_active_vrpred ? _T_2242 & _T_7 | ~_T_7 & _T_3682 : _T_3682;	// sequencer-master.scala:131:52, :183:52
      wire _T_3691 = io_op_bits_active_vrpred ? _T_2246 & _T_7 | ~_T_7 & _T_3683 : _T_3683;	// sequencer-master.scala:131:52, :183:52
      wire _T_3692 = io_op_bits_active_vrpred ? _T_2250 & _T_7 | ~_T_7 & _T_3684 : _T_3684;	// sequencer-master.scala:131:52, :183:52
      wire _T_3693 = io_op_bits_active_vrpred ? _T_2254 & _T_7 | ~_T_7 & _T_3685 : _T_3685;	// sequencer-master.scala:131:52, :183:52
      wire _T_3694 = io_op_bits_active_vrpred ? _T_2258 & _T_7 | ~_T_7 & _T_3686 : _T_3686;	// sequencer-master.scala:131:52, :183:52
      wire _T_3695 = io_op_bits_active_vrpred ? _T_2262 & _T_7 | ~_T_7 & _T_3687 : _T_3687;	// sequencer-master.scala:131:52, :183:52
      wire _T_3696 = io_op_bits_active_vrpred ? _T_2266 & _T_7 | ~_T_7 & _T_3688 : _T_3688;	// sequencer-master.scala:131:52, :183:52
      wire _T_3697 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_7 | ~_T_7 & _T_3665 : _T_3665);	// sequencer-master.scala:132:52, :184:52
      wire _T_3698 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_7 | ~_T_7 & _T_3673 : _T_3673);	// sequencer-master.scala:133:52, :185:52
      wire _T_3699 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_7 | ~_T_7 & _T_3666 : _T_3666);	// sequencer-master.scala:132:52, :184:52
      wire _T_3700 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_7 | ~_T_7 & _T_3674 : _T_3674);	// sequencer-master.scala:133:52, :185:52
      wire _T_3701 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_7 | ~_T_7 & _T_3667 : _T_3667);	// sequencer-master.scala:132:52, :184:52
      wire _T_3702 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_7 | ~_T_7 & _T_3675 : _T_3675);	// sequencer-master.scala:133:52, :185:52
      wire _T_3703 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_7 | ~_T_7 & _T_3668 : _T_3668);	// sequencer-master.scala:132:52, :184:52
      wire _T_3704 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_7 | ~_T_7 & _T_3676 : _T_3676);	// sequencer-master.scala:133:52, :185:52
      wire _T_3705 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_7 | ~_T_7 & _T_3669 : _T_3669);	// sequencer-master.scala:132:52, :184:52
      wire _T_3706 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_7 | ~_T_7 & _T_3677 : _T_3677);	// sequencer-master.scala:133:52, :185:52
      wire _T_3707 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_7 | ~_T_7 & _T_3670 : _T_3670);	// sequencer-master.scala:132:52, :184:52
      wire _T_3708 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_7 | ~_T_7 & _T_3678 : _T_3678);	// sequencer-master.scala:133:52, :185:52
      wire _T_3709 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_7 | ~_T_7 & _T_3671 : _T_3671);	// sequencer-master.scala:132:52, :184:52
      wire _T_3710 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_7 | ~_T_7 & _T_3679 : _T_3679);	// sequencer-master.scala:133:52, :185:52
      wire _T_3711 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_7 | ~_T_7 & _T_3672 : _T_3672);	// sequencer-master.scala:132:52, :184:52
      wire _T_3712 = (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_7 | ~_T_7 & _T_3680 : _T_3680);	// sequencer-master.scala:133:52, :185:52
      wire _T_3713 = io_op_bits_active_vrfirst ? _T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 & _T_3689 : _T_3689;	// sequencer-master.scala:131:52, :183:52
      wire _T_3714 = io_op_bits_active_vrfirst ? _T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 & _T_3690 : _T_3690;	// sequencer-master.scala:131:52, :183:52
      wire _T_3715 = io_op_bits_active_vrfirst ? _T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 & _T_3691 : _T_3691;	// sequencer-master.scala:131:52, :183:52
      wire _T_3716 = io_op_bits_active_vrfirst ? _T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 & _T_3692 : _T_3692;	// sequencer-master.scala:131:52, :183:52
      wire _T_3717 = io_op_bits_active_vrfirst ? _T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 & _T_3693 : _T_3693;	// sequencer-master.scala:131:52, :183:52
      wire _T_3718 = io_op_bits_active_vrfirst ? _T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 & _T_3694 : _T_3694;	// sequencer-master.scala:131:52, :183:52
      wire _T_3719 = io_op_bits_active_vrfirst ? _T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 & _T_3695 : _T_3695;	// sequencer-master.scala:131:52, :183:52
      wire _T_3720 = io_op_bits_active_vrfirst ? _T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 & _T_3696 : _T_3696;	// sequencer-master.scala:131:52, :183:52
      wire _T_3721 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_132 | _T_2279 & _T_294 | _T_2238 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2269 & _T_7 | _T_2238 & _T_7 | ~_T_7 & _T_3713)) : _T_3713;	// sequencer-master.scala:131:52, :183:52
      wire _T_3722 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_133 | _T_2280 & _T_294 | _T_2242 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2270 & _T_7 | _T_2242 & _T_7 | ~_T_7 & _T_3714)) : _T_3714;	// sequencer-master.scala:131:52, :183:52
      wire _T_3723 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_134 | _T_2281 & _T_294 | _T_2246 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2271 & _T_7 | _T_2246 & _T_7 | ~_T_7 & _T_3715)) : _T_3715;	// sequencer-master.scala:131:52, :183:52
      wire _T_3724 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_135 | _T_2282 & _T_294 | _T_2250 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2272 & _T_7 | _T_2250 & _T_7 | ~_T_7 & _T_3716)) : _T_3716;	// sequencer-master.scala:131:52, :183:52
      wire _T_3725 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_136 | _T_2283 & _T_294 | _T_2254 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2273 & _T_7 | _T_2254 & _T_7 | ~_T_7 & _T_3717)) : _T_3717;	// sequencer-master.scala:131:52, :183:52
      wire _T_3726 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_137 | _T_2284 & _T_294 | _T_2258 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2274 & _T_7 | _T_2258 & _T_7 | ~_T_7 & _T_3718)) : _T_3718;	// sequencer-master.scala:131:52, :183:52
      wire _T_3727 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & _T_138 | _T_2285 & _T_294 | _T_2262 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2275 & _T_7 | _T_2262 & _T_7 | ~_T_7 & _T_3719)) : _T_3719;	// sequencer-master.scala:131:52, :183:52
      wire _T_3728 = io_op_bits_active_vamo ? ~_T_317 & (_T_294 & &_T_0 | _T_2286 & _T_294 | _T_2266 & _T_294 |
                ~_T_294 & ~_T_135 & (_T_2276 & _T_7 | _T_2266 & _T_7 | ~_T_7 & _T_3720)) : _T_3720;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3729 = io_op_bits_active_vamo ? _T_2308 & _T_317 | ~_T_317 & ~_T_294 & (_T_2308 & _T_135 | ~_T_135
                & ~_T_7 & _T_3697) : _T_3697;	// sequencer-master.scala:132:52, :184:52
      wire _T_3730 = io_op_bits_active_vamo ? _T_2309 & _T_317 | ~_T_317 & ~_T_294 & (_T_2309 & _T_135 | ~_T_135
                & ~_T_7 & _T_3699) : _T_3699;	// sequencer-master.scala:132:52, :184:52
      wire _T_3731 = io_op_bits_active_vamo ? _T_2310 & _T_317 | ~_T_317 & ~_T_294 & (_T_2310 & _T_135 | ~_T_135
                & ~_T_7 & _T_3701) : _T_3701;	// sequencer-master.scala:132:52, :184:52
      wire _T_3732 = io_op_bits_active_vamo ? _T_2311 & _T_317 | ~_T_317 & ~_T_294 & (_T_2311 & _T_135 | ~_T_135
                & ~_T_7 & _T_3703) : _T_3703;	// sequencer-master.scala:132:52, :184:52
      wire _T_3733 = io_op_bits_active_vamo ? _T_2312 & _T_317 | ~_T_317 & ~_T_294 & (_T_2312 & _T_135 | ~_T_135
                & ~_T_7 & _T_3705) : _T_3705;	// sequencer-master.scala:132:52, :184:52
      wire _T_3734 = io_op_bits_active_vamo ? _T_2313 & _T_317 | ~_T_317 & ~_T_294 & (_T_2313 & _T_135 | ~_T_135
                & ~_T_7 & _T_3707) : _T_3707;	// sequencer-master.scala:132:52, :184:52
      wire _T_3735 = io_op_bits_active_vamo ? _T_2314 & _T_317 | ~_T_317 & ~_T_294 & (_T_2314 & _T_135 | ~_T_135
                & ~_T_7 & _T_3709) : _T_3709;	// sequencer-master.scala:132:52, :184:52
      wire _T_3736 = io_op_bits_active_vamo ? _T_2315 & _T_317 | ~_T_317 & ~_T_294 & (_T_2315 & _T_135 | ~_T_135
                & ~_T_7 & _T_3711) : _T_3711;	// sequencer-master.scala:132:52, :184:52
      wire _T_3737 = io_op_bits_active_vamo ? _T_2299 & _T_317 | ~_T_317 & ~_T_294 & (_T_2299 & _T_135 | ~_T_135
                & ~_T_7 & _T_3698) : _T_3698;	// sequencer-master.scala:133:52, :185:52
      wire _T_3738 = io_op_bits_active_vamo ? _T_2300 & _T_317 | ~_T_317 & ~_T_294 & (_T_2300 & _T_135 | ~_T_135
                & ~_T_7 & _T_3700) : _T_3700;	// sequencer-master.scala:133:52, :185:52
      wire _T_3739 = io_op_bits_active_vamo ? _T_2301 & _T_317 | ~_T_317 & ~_T_294 & (_T_2301 & _T_135 | ~_T_135
                & ~_T_7 & _T_3702) : _T_3702;	// sequencer-master.scala:133:52, :185:52
      wire _T_3740 = io_op_bits_active_vamo ? _T_2302 & _T_317 | ~_T_317 & ~_T_294 & (_T_2302 & _T_135 | ~_T_135
                & ~_T_7 & _T_3704) : _T_3704;	// sequencer-master.scala:133:52, :185:52
      wire _T_3741 = io_op_bits_active_vamo ? _T_2303 & _T_317 | ~_T_317 & ~_T_294 & (_T_2303 & _T_135 | ~_T_135
                & ~_T_7 & _T_3706) : _T_3706;	// sequencer-master.scala:133:52, :185:52
      wire _T_3742 = io_op_bits_active_vamo ? _T_2304 & _T_317 | ~_T_317 & ~_T_294 & (_T_2304 & _T_135 | ~_T_135
                & ~_T_7 & _T_3708) : _T_3708;	// sequencer-master.scala:133:52, :185:52
      wire _T_3743 = io_op_bits_active_vamo ? _T_2305 & _T_317 | ~_T_317 & ~_T_294 & (_T_2305 & _T_135 | ~_T_135
                & ~_T_7 & _T_3710) : _T_3710;	// sequencer-master.scala:133:52, :185:52
      wire _T_3744 = io_op_bits_active_vamo ? _T_2306 & _T_317 | ~_T_317 & ~_T_294 & (_T_2306 & _T_135 | ~_T_135
                & ~_T_7 & _T_3712) : _T_3712;	// sequencer-master.scala:133:52, :185:52
      wire _T_3745 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2279 & _T_7 | _T_2238 & _T_7 | ~_T_7 &
                _T_3721) : _T_3721;	// sequencer-master.scala:131:52, :183:52
      wire _T_3746 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2280 & _T_7 | _T_2242 & _T_7 | ~_T_7 &
                _T_3722) : _T_3722;	// sequencer-master.scala:131:52, :183:52
      wire _T_3747 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2281 & _T_7 | _T_2246 & _T_7 | ~_T_7 &
                _T_3723) : _T_3723;	// sequencer-master.scala:131:52, :183:52
      wire _T_3748 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2282 & _T_7 | _T_2250 & _T_7 | ~_T_7 &
                _T_3724) : _T_3724;	// sequencer-master.scala:131:52, :183:52
      wire _T_3749 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2283 & _T_7 | _T_2254 & _T_7 | ~_T_7 &
                _T_3725) : _T_3725;	// sequencer-master.scala:131:52, :183:52
      wire _T_3750 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2284 & _T_7 | _T_2258 & _T_7 | ~_T_7 &
                _T_3726) : _T_3726;	// sequencer-master.scala:131:52, :183:52
      wire _T_3751 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2285 & _T_7 | _T_2262 & _T_7 | ~_T_7 &
                _T_3727) : _T_3727;	// sequencer-master.scala:131:52, :183:52
      wire _T_3752 = io_op_bits_active_vldx ? ~_T_294 & ~_T_135 & (_T_2286 & _T_7 | _T_2266 & _T_7 | ~_T_7 &
                _T_3728) : _T_3728;	// sequencer-master.scala:131:52, :183:52
      wire _T_3753 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2308 &
                _T_294 | ~_T_294 & (_T_2308 & _T_135 | ~_T_135 & ~_T_7 & _T_3729) : _T_3729);	// sequencer-master.scala:132:52, :184:52
      wire _T_3754 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2299 &
                _T_294 | ~_T_294 & (_T_2299 & _T_135 | ~_T_135 & ~_T_7 & _T_3737) : _T_3737);	// sequencer-master.scala:133:52, :185:52
      wire _T_3755 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2309 &
                _T_294 | ~_T_294 & (_T_2309 & _T_135 | ~_T_135 & ~_T_7 & _T_3730) : _T_3730);	// sequencer-master.scala:132:52, :184:52
      wire _T_3756 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2300 &
                _T_294 | ~_T_294 & (_T_2300 & _T_135 | ~_T_135 & ~_T_7 & _T_3738) : _T_3738);	// sequencer-master.scala:133:52, :185:52
      wire _T_3757 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2310 &
                _T_294 | ~_T_294 & (_T_2310 & _T_135 | ~_T_135 & ~_T_7 & _T_3731) : _T_3731);	// sequencer-master.scala:132:52, :184:52
      wire _T_3758 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2301 &
                _T_294 | ~_T_294 & (_T_2301 & _T_135 | ~_T_135 & ~_T_7 & _T_3739) : _T_3739);	// sequencer-master.scala:133:52, :185:52
      wire _T_3759 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2311 &
                _T_294 | ~_T_294 & (_T_2311 & _T_135 | ~_T_135 & ~_T_7 & _T_3732) : _T_3732);	// sequencer-master.scala:132:52, :184:52
      wire _T_3760 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2302 &
                _T_294 | ~_T_294 & (_T_2302 & _T_135 | ~_T_135 & ~_T_7 & _T_3740) : _T_3740);	// sequencer-master.scala:133:52, :185:52
      wire _T_3761 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2312 &
                _T_294 | ~_T_294 & (_T_2312 & _T_135 | ~_T_135 & ~_T_7 & _T_3733) : _T_3733);	// sequencer-master.scala:132:52, :184:52
      wire _T_3762 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2303 &
                _T_294 | ~_T_294 & (_T_2303 & _T_135 | ~_T_135 & ~_T_7 & _T_3741) : _T_3741);	// sequencer-master.scala:133:52, :185:52
      wire _T_3763 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2313 &
                _T_294 | ~_T_294 & (_T_2313 & _T_135 | ~_T_135 & ~_T_7 & _T_3734) : _T_3734);	// sequencer-master.scala:132:52, :184:52
      wire _T_3764 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2304 &
                _T_294 | ~_T_294 & (_T_2304 & _T_135 | ~_T_135 & ~_T_7 & _T_3742) : _T_3742);	// sequencer-master.scala:133:52, :185:52
      wire _T_3765 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2314 &
                _T_294 | ~_T_294 & (_T_2314 & _T_135 | ~_T_135 & ~_T_7 & _T_3735) : _T_3735);	// sequencer-master.scala:132:52, :184:52
      wire _T_3766 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2305 &
                _T_294 | ~_T_294 & (_T_2305 & _T_135 | ~_T_135 & ~_T_7 & _T_3743) : _T_3743);	// sequencer-master.scala:133:52, :185:52
      wire _T_3767 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2315 &
                _T_294 | ~_T_294 & (_T_2315 & _T_135 | ~_T_135 & ~_T_7 & _T_3736) : _T_3736);	// sequencer-master.scala:132:52, :184:52
      wire _T_3768 = (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vldx ? _T_2306 &
                _T_294 | ~_T_294 & (_T_2306 & _T_135 | ~_T_135 & ~_T_7 & _T_3744) : _T_3744);	// sequencer-master.scala:133:52, :185:52
      wire _T_3769 = io_op_bits_active_vstx ? _T_294 & _T_132 | _T_2299 & _T_294 | _T_2238 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2279 & _T_7 | _T_2238 & _T_7 | ~_T_7 & _T_3745) : _T_3745;	// sequencer-master.scala:131:52, :183:52
      wire _T_3770 = io_op_bits_active_vstx ? _T_294 & _T_133 | _T_2300 & _T_294 | _T_2242 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2280 & _T_7 | _T_2242 & _T_7 | ~_T_7 & _T_3746) : _T_3746;	// sequencer-master.scala:131:52, :183:52
      wire _T_3771 = io_op_bits_active_vstx ? _T_294 & _T_134 | _T_2301 & _T_294 | _T_2246 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2281 & _T_7 | _T_2246 & _T_7 | ~_T_7 & _T_3747) : _T_3747;	// sequencer-master.scala:131:52, :183:52
      wire _T_3772 = io_op_bits_active_vstx ? _T_294 & _T_135 | _T_2302 & _T_294 | _T_2250 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2282 & _T_7 | _T_2250 & _T_7 | ~_T_7 & _T_3748) : _T_3748;	// sequencer-master.scala:131:52, :183:52
      wire _T_3773 = io_op_bits_active_vstx ? _T_294 & _T_136 | _T_2303 & _T_294 | _T_2254 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2283 & _T_7 | _T_2254 & _T_7 | ~_T_7 & _T_3749) : _T_3749;	// sequencer-master.scala:131:52, :183:52
      wire _T_3774 = io_op_bits_active_vstx ? _T_294 & _T_137 | _T_2304 & _T_294 | _T_2258 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2284 & _T_7 | _T_2258 & _T_7 | ~_T_7 & _T_3750) : _T_3750;	// sequencer-master.scala:131:52, :183:52
      wire _T_3775 = io_op_bits_active_vstx ? _T_294 & _T_138 | _T_2305 & _T_294 | _T_2262 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2285 & _T_7 | _T_2262 & _T_7 | ~_T_7 & _T_3751) : _T_3751;	// sequencer-master.scala:131:52, :183:52
      wire _T_3776 = io_op_bits_active_vstx ? _T_294 & &_T_0 | _T_2306 & _T_294 | _T_2266 & _T_294 | ~_T_294 &
                ~_T_135 & (_T_2286 & _T_7 | _T_2266 & _T_7 | ~_T_7 & _T_3752) : _T_3752;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_3777 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2238 & _T_7 | ~_T_7 & _T_3769) : _T_3769;	// sequencer-master.scala:131:52, :183:52
      wire _T_3778 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2242 & _T_7 | ~_T_7 & _T_3770) : _T_3770;	// sequencer-master.scala:131:52, :183:52
      wire _T_3779 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2246 & _T_7 | ~_T_7 & _T_3771) : _T_3771;	// sequencer-master.scala:131:52, :183:52
      wire _T_3780 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2250 & _T_7 | ~_T_7 & _T_3772) : _T_3772;	// sequencer-master.scala:131:52, :183:52
      wire _T_3781 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2254 & _T_7 | ~_T_7 & _T_3773) : _T_3773;	// sequencer-master.scala:131:52, :183:52
      wire _T_3782 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2258 & _T_7 | ~_T_7 & _T_3774) : _T_3774;	// sequencer-master.scala:131:52, :183:52
      wire _T_3783 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2262 & _T_7 | ~_T_7 & _T_3775) : _T_3775;	// sequencer-master.scala:131:52, :183:52
      wire _T_3784 = io_op_bits_active_vld ? ~_T_294 & ~_T_135 & (_T_2266 & _T_7 | ~_T_7 & _T_3776) : _T_3776;	// sequencer-master.scala:131:52, :183:52
      wire _T_3785 = io_op_bits_active_vint ? _T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 &
                e_4_raw_0 : e_4_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_3786 = io_op_bits_active_vint ? _T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 &
                e_4_raw_1 : e_4_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_3787 = io_op_bits_active_vint ? _T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 &
                e_4_raw_2 : e_4_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_3788 = io_op_bits_active_vint ? _T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 &
                e_4_raw_3 : e_4_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_3789 = io_op_bits_active_vint ? _T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 &
                e_4_raw_4 : e_4_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_3790 = io_op_bits_active_vint ? _T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 &
                e_4_raw_5 : e_4_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_3791 = io_op_bits_active_vint ? _T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 &
                e_4_raw_6 : e_4_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_3792 = io_op_bits_active_vint ? _T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 &
                e_4_raw_7 : e_4_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_3793 = io_op_bits_active_vint ? _T_2308 & _T_8 | ~_T_8 & e_4_war_0 : e_4_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_3794 = io_op_bits_active_vint ? _T_2309 & _T_8 | ~_T_8 & e_4_war_1 : e_4_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_3795 = io_op_bits_active_vint ? _T_2310 & _T_8 | ~_T_8 & e_4_war_2 : e_4_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_3796 = io_op_bits_active_vint ? _T_2311 & _T_8 | ~_T_8 & e_4_war_3 : e_4_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_3797 = io_op_bits_active_vint ? _T_2312 & _T_8 | ~_T_8 & e_4_war_4 : e_4_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_3798 = io_op_bits_active_vint ? _T_2313 & _T_8 | ~_T_8 & e_4_war_5 : e_4_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_3799 = io_op_bits_active_vint ? _T_2314 & _T_8 | ~_T_8 & e_4_war_6 : e_4_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_3800 = io_op_bits_active_vint ? _T_2315 & _T_8 | ~_T_8 & e_4_war_7 : e_4_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_3801 = io_op_bits_active_vint ? _T_2299 & _T_8 | ~_T_8 & e_4_waw_0 : e_4_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_3802 = io_op_bits_active_vint ? _T_2300 & _T_8 | ~_T_8 & e_4_waw_1 : e_4_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_3803 = io_op_bits_active_vint ? _T_2301 & _T_8 | ~_T_8 & e_4_waw_2 : e_4_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_3804 = io_op_bits_active_vint ? _T_2302 & _T_8 | ~_T_8 & e_4_waw_3 : e_4_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_3805 = io_op_bits_active_vint ? _T_2303 & _T_8 | ~_T_8 & e_4_waw_4 : e_4_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_3806 = io_op_bits_active_vint ? _T_2304 & _T_8 | ~_T_8 & e_4_waw_5 : e_4_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_3807 = io_op_bits_active_vint ? _T_2305 & _T_8 | ~_T_8 & e_4_waw_6 : e_4_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_3808 = io_op_bits_active_vint ? _T_2306 & _T_8 | ~_T_8 & e_4_waw_7 : e_4_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_3809 = io_op_bits_active_vipred ? _T_2289 & _T_8 | _T_2279 & _T_8 | _T_2269 & _T_8 | ~_T_8 &
                _T_3785 : _T_3785;	// sequencer-master.scala:131:52, :183:52
      wire _T_3810 = io_op_bits_active_vipred ? _T_2290 & _T_8 | _T_2280 & _T_8 | _T_2270 & _T_8 | ~_T_8 &
                _T_3786 : _T_3786;	// sequencer-master.scala:131:52, :183:52
      wire _T_3811 = io_op_bits_active_vipred ? _T_2291 & _T_8 | _T_2281 & _T_8 | _T_2271 & _T_8 | ~_T_8 &
                _T_3787 : _T_3787;	// sequencer-master.scala:131:52, :183:52
      wire _T_3812 = io_op_bits_active_vipred ? _T_2292 & _T_8 | _T_2282 & _T_8 | _T_2272 & _T_8 | ~_T_8 &
                _T_3788 : _T_3788;	// sequencer-master.scala:131:52, :183:52
      wire _T_3813 = io_op_bits_active_vipred ? _T_2293 & _T_8 | _T_2283 & _T_8 | _T_2273 & _T_8 | ~_T_8 &
                _T_3789 : _T_3789;	// sequencer-master.scala:131:52, :183:52
      wire _T_3814 = io_op_bits_active_vipred ? _T_2294 & _T_8 | _T_2284 & _T_8 | _T_2274 & _T_8 | ~_T_8 &
                _T_3790 : _T_3790;	// sequencer-master.scala:131:52, :183:52
      wire _T_3815 = io_op_bits_active_vipred ? _T_2295 & _T_8 | _T_2285 & _T_8 | _T_2275 & _T_8 | ~_T_8 &
                _T_3791 : _T_3791;	// sequencer-master.scala:131:52, :183:52
      wire _T_3816 = io_op_bits_active_vipred ? _T_2296 & _T_8 | _T_2286 & _T_8 | _T_2276 & _T_8 | ~_T_8 &
                _T_3792 : _T_3792;	// sequencer-master.scala:131:52, :183:52
      wire _T_3817 = io_op_bits_active_vipred ? _T_2308 & _T_8 | ~_T_8 & _T_3793 : _T_3793;	// sequencer-master.scala:132:52, :184:52
      wire _T_3818 = io_op_bits_active_vipred ? _T_2309 & _T_8 | ~_T_8 & _T_3794 : _T_3794;	// sequencer-master.scala:132:52, :184:52
      wire _T_3819 = io_op_bits_active_vipred ? _T_2310 & _T_8 | ~_T_8 & _T_3795 : _T_3795;	// sequencer-master.scala:132:52, :184:52
      wire _T_3820 = io_op_bits_active_vipred ? _T_2311 & _T_8 | ~_T_8 & _T_3796 : _T_3796;	// sequencer-master.scala:132:52, :184:52
      wire _T_3821 = io_op_bits_active_vipred ? _T_2312 & _T_8 | ~_T_8 & _T_3797 : _T_3797;	// sequencer-master.scala:132:52, :184:52
      wire _T_3822 = io_op_bits_active_vipred ? _T_2313 & _T_8 | ~_T_8 & _T_3798 : _T_3798;	// sequencer-master.scala:132:52, :184:52
      wire _T_3823 = io_op_bits_active_vipred ? _T_2314 & _T_8 | ~_T_8 & _T_3799 : _T_3799;	// sequencer-master.scala:132:52, :184:52
      wire _T_3824 = io_op_bits_active_vipred ? _T_2315 & _T_8 | ~_T_8 & _T_3800 : _T_3800;	// sequencer-master.scala:132:52, :184:52
      wire _T_3825 = io_op_bits_active_vipred ? _T_2299 & _T_8 | ~_T_8 & _T_3801 : _T_3801;	// sequencer-master.scala:133:52, :185:52
      wire _T_3826 = io_op_bits_active_vipred ? _T_2300 & _T_8 | ~_T_8 & _T_3802 : _T_3802;	// sequencer-master.scala:133:52, :185:52
      wire _T_3827 = io_op_bits_active_vipred ? _T_2301 & _T_8 | ~_T_8 & _T_3803 : _T_3803;	// sequencer-master.scala:133:52, :185:52
      wire _T_3828 = io_op_bits_active_vipred ? _T_2302 & _T_8 | ~_T_8 & _T_3804 : _T_3804;	// sequencer-master.scala:133:52, :185:52
      wire _T_3829 = io_op_bits_active_vipred ? _T_2303 & _T_8 | ~_T_8 & _T_3805 : _T_3805;	// sequencer-master.scala:133:52, :185:52
      wire _T_3830 = io_op_bits_active_vipred ? _T_2304 & _T_8 | ~_T_8 & _T_3806 : _T_3806;	// sequencer-master.scala:133:52, :185:52
      wire _T_3831 = io_op_bits_active_vipred ? _T_2305 & _T_8 | ~_T_8 & _T_3807 : _T_3807;	// sequencer-master.scala:133:52, :185:52
      wire _T_3832 = io_op_bits_active_vipred ? _T_2306 & _T_8 | ~_T_8 & _T_3808 : _T_3808;	// sequencer-master.scala:133:52, :185:52
      wire _T_3833 = io_op_bits_active_vimul ? _T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 &
                _T_3809 : _T_3809;	// sequencer-master.scala:131:52, :183:52
      wire _T_3834 = io_op_bits_active_vimul ? _T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 &
                _T_3810 : _T_3810;	// sequencer-master.scala:131:52, :183:52
      wire _T_3835 = io_op_bits_active_vimul ? _T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 &
                _T_3811 : _T_3811;	// sequencer-master.scala:131:52, :183:52
      wire _T_3836 = io_op_bits_active_vimul ? _T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 &
                _T_3812 : _T_3812;	// sequencer-master.scala:131:52, :183:52
      wire _T_3837 = io_op_bits_active_vimul ? _T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 &
                _T_3813 : _T_3813;	// sequencer-master.scala:131:52, :183:52
      wire _T_3838 = io_op_bits_active_vimul ? _T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 &
                _T_3814 : _T_3814;	// sequencer-master.scala:131:52, :183:52
      wire _T_3839 = io_op_bits_active_vimul ? _T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 &
                _T_3815 : _T_3815;	// sequencer-master.scala:131:52, :183:52
      wire _T_3840 = io_op_bits_active_vimul ? _T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 &
                _T_3816 : _T_3816;	// sequencer-master.scala:131:52, :183:52
      wire _T_3841 = io_op_bits_active_vimul ? _T_2308 & _T_8 | ~_T_8 & _T_3817 : _T_3817;	// sequencer-master.scala:132:52, :184:52
      wire _T_3842 = io_op_bits_active_vimul ? _T_2309 & _T_8 | ~_T_8 & _T_3818 : _T_3818;	// sequencer-master.scala:132:52, :184:52
      wire _T_3843 = io_op_bits_active_vimul ? _T_2310 & _T_8 | ~_T_8 & _T_3819 : _T_3819;	// sequencer-master.scala:132:52, :184:52
      wire _T_3844 = io_op_bits_active_vimul ? _T_2311 & _T_8 | ~_T_8 & _T_3820 : _T_3820;	// sequencer-master.scala:132:52, :184:52
      wire _T_3845 = io_op_bits_active_vimul ? _T_2312 & _T_8 | ~_T_8 & _T_3821 : _T_3821;	// sequencer-master.scala:132:52, :184:52
      wire _T_3846 = io_op_bits_active_vimul ? _T_2313 & _T_8 | ~_T_8 & _T_3822 : _T_3822;	// sequencer-master.scala:132:52, :184:52
      wire _T_3847 = io_op_bits_active_vimul ? _T_2314 & _T_8 | ~_T_8 & _T_3823 : _T_3823;	// sequencer-master.scala:132:52, :184:52
      wire _T_3848 = io_op_bits_active_vimul ? _T_2315 & _T_8 | ~_T_8 & _T_3824 : _T_3824;	// sequencer-master.scala:132:52, :184:52
      wire _T_3849 = io_op_bits_active_vimul ? _T_2299 & _T_8 | ~_T_8 & _T_3825 : _T_3825;	// sequencer-master.scala:133:52, :185:52
      wire _T_3850 = io_op_bits_active_vimul ? _T_2300 & _T_8 | ~_T_8 & _T_3826 : _T_3826;	// sequencer-master.scala:133:52, :185:52
      wire _T_3851 = io_op_bits_active_vimul ? _T_2301 & _T_8 | ~_T_8 & _T_3827 : _T_3827;	// sequencer-master.scala:133:52, :185:52
      wire _T_3852 = io_op_bits_active_vimul ? _T_2302 & _T_8 | ~_T_8 & _T_3828 : _T_3828;	// sequencer-master.scala:133:52, :185:52
      wire _T_3853 = io_op_bits_active_vimul ? _T_2303 & _T_8 | ~_T_8 & _T_3829 : _T_3829;	// sequencer-master.scala:133:52, :185:52
      wire _T_3854 = io_op_bits_active_vimul ? _T_2304 & _T_8 | ~_T_8 & _T_3830 : _T_3830;	// sequencer-master.scala:133:52, :185:52
      wire _T_3855 = io_op_bits_active_vimul ? _T_2305 & _T_8 | ~_T_8 & _T_3831 : _T_3831;	// sequencer-master.scala:133:52, :185:52
      wire _T_3856 = io_op_bits_active_vimul ? _T_2306 & _T_8 | ~_T_8 & _T_3832 : _T_3832;	// sequencer-master.scala:133:52, :185:52
      wire _T_3857 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8 |
                ~_T_8 & _T_3833) : _T_3833;	// sequencer-master.scala:131:52, :183:52
      wire _T_3858 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8 |
                ~_T_8 & _T_3834) : _T_3834;	// sequencer-master.scala:131:52, :183:52
      wire _T_3859 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8 |
                ~_T_8 & _T_3835) : _T_3835;	// sequencer-master.scala:131:52, :183:52
      wire _T_3860 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8 |
                ~_T_8 & _T_3836) : _T_3836;	// sequencer-master.scala:131:52, :183:52
      wire _T_3861 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8 |
                ~_T_8 & _T_3837) : _T_3837;	// sequencer-master.scala:131:52, :183:52
      wire _T_3862 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8 |
                ~_T_8 & _T_3838) : _T_3838;	// sequencer-master.scala:131:52, :183:52
      wire _T_3863 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8 |
                ~_T_8 & _T_3839) : _T_3839;	// sequencer-master.scala:131:52, :183:52
      wire _T_3864 = io_op_bits_active_vidiv ? ~_T_136 & (_T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8 |
                ~_T_8 & _T_3840) : _T_3840;	// sequencer-master.scala:131:52, :183:52
      wire _T_3865 = io_op_bits_active_vidiv ? _T_2308 & _T_136 | ~_T_136 & (_T_2308 & _T_8 | ~_T_8 & _T_3841) :
                _T_3841;	// sequencer-master.scala:132:52, :184:52
      wire _T_3866 = io_op_bits_active_vidiv ? _T_2309 & _T_136 | ~_T_136 & (_T_2309 & _T_8 | ~_T_8 & _T_3842) :
                _T_3842;	// sequencer-master.scala:132:52, :184:52
      wire _T_3867 = io_op_bits_active_vidiv ? _T_2310 & _T_136 | ~_T_136 & (_T_2310 & _T_8 | ~_T_8 & _T_3843) :
                _T_3843;	// sequencer-master.scala:132:52, :184:52
      wire _T_3868 = io_op_bits_active_vidiv ? _T_2311 & _T_136 | ~_T_136 & (_T_2311 & _T_8 | ~_T_8 & _T_3844) :
                _T_3844;	// sequencer-master.scala:132:52, :184:52
      wire _T_3869 = io_op_bits_active_vidiv ? _T_2312 & _T_136 | ~_T_136 & (_T_2312 & _T_8 | ~_T_8 & _T_3845) :
                _T_3845;	// sequencer-master.scala:132:52, :184:52
      wire _T_3870 = io_op_bits_active_vidiv ? _T_2313 & _T_136 | ~_T_136 & (_T_2313 & _T_8 | ~_T_8 & _T_3846) :
                _T_3846;	// sequencer-master.scala:132:52, :184:52
      wire _T_3871 = io_op_bits_active_vidiv ? _T_2314 & _T_136 | ~_T_136 & (_T_2314 & _T_8 | ~_T_8 & _T_3847) :
                _T_3847;	// sequencer-master.scala:132:52, :184:52
      wire _T_3872 = io_op_bits_active_vidiv ? _T_2315 & _T_136 | ~_T_136 & (_T_2315 & _T_8 | ~_T_8 & _T_3848) :
                _T_3848;	// sequencer-master.scala:132:52, :184:52
      wire _T_3873 = io_op_bits_active_vidiv ? _T_2299 & _T_136 | ~_T_136 & (_T_2299 & _T_8 | ~_T_8 & _T_3849) :
                _T_3849;	// sequencer-master.scala:133:52, :185:52
      wire _T_3874 = io_op_bits_active_vidiv ? _T_2300 & _T_136 | ~_T_136 & (_T_2300 & _T_8 | ~_T_8 & _T_3850) :
                _T_3850;	// sequencer-master.scala:133:52, :185:52
      wire _T_3875 = io_op_bits_active_vidiv ? _T_2301 & _T_136 | ~_T_136 & (_T_2301 & _T_8 | ~_T_8 & _T_3851) :
                _T_3851;	// sequencer-master.scala:133:52, :185:52
      wire _T_3876 = io_op_bits_active_vidiv ? _T_2302 & _T_136 | ~_T_136 & (_T_2302 & _T_8 | ~_T_8 & _T_3852) :
                _T_3852;	// sequencer-master.scala:133:52, :185:52
      wire _T_3877 = io_op_bits_active_vidiv ? _T_2303 & _T_136 | ~_T_136 & (_T_2303 & _T_8 | ~_T_8 & _T_3853) :
                _T_3853;	// sequencer-master.scala:133:52, :185:52
      wire _T_3878 = io_op_bits_active_vidiv ? _T_2304 & _T_136 | ~_T_136 & (_T_2304 & _T_8 | ~_T_8 & _T_3854) :
                _T_3854;	// sequencer-master.scala:133:52, :185:52
      wire _T_3879 = io_op_bits_active_vidiv ? _T_2305 & _T_136 | ~_T_136 & (_T_2305 & _T_8 | ~_T_8 & _T_3855) :
                _T_3855;	// sequencer-master.scala:133:52, :185:52
      wire _T_3880 = io_op_bits_active_vidiv ? _T_2306 & _T_136 | ~_T_136 & (_T_2306 & _T_8 | ~_T_8 & _T_3856) :
                _T_3856;	// sequencer-master.scala:133:52, :185:52
      wire _T_3881 = io_op_bits_active_vfma ? _T_2289 & _T_8 | _T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8
                | ~_T_8 & _T_3857 : _T_3857;	// sequencer-master.scala:131:52, :183:52
      wire _T_3882 = io_op_bits_active_vfma ? _T_2290 & _T_8 | _T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8
                | ~_T_8 & _T_3858 : _T_3858;	// sequencer-master.scala:131:52, :183:52
      wire _T_3883 = io_op_bits_active_vfma ? _T_2291 & _T_8 | _T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8
                | ~_T_8 & _T_3859 : _T_3859;	// sequencer-master.scala:131:52, :183:52
      wire _T_3884 = io_op_bits_active_vfma ? _T_2292 & _T_8 | _T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8
                | ~_T_8 & _T_3860 : _T_3860;	// sequencer-master.scala:131:52, :183:52
      wire _T_3885 = io_op_bits_active_vfma ? _T_2293 & _T_8 | _T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8
                | ~_T_8 & _T_3861 : _T_3861;	// sequencer-master.scala:131:52, :183:52
      wire _T_3886 = io_op_bits_active_vfma ? _T_2294 & _T_8 | _T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8
                | ~_T_8 & _T_3862 : _T_3862;	// sequencer-master.scala:131:52, :183:52
      wire _T_3887 = io_op_bits_active_vfma ? _T_2295 & _T_8 | _T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8
                | ~_T_8 & _T_3863 : _T_3863;	// sequencer-master.scala:131:52, :183:52
      wire _T_3888 = io_op_bits_active_vfma ? _T_2296 & _T_8 | _T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8
                | ~_T_8 & _T_3864 : _T_3864;	// sequencer-master.scala:131:52, :183:52
      wire _T_3889 = io_op_bits_active_vfma ? _T_2308 & _T_8 | ~_T_8 & _T_3865 : _T_3865;	// sequencer-master.scala:132:52, :184:52
      wire _T_3890 = io_op_bits_active_vfma ? _T_2309 & _T_8 | ~_T_8 & _T_3866 : _T_3866;	// sequencer-master.scala:132:52, :184:52
      wire _T_3891 = io_op_bits_active_vfma ? _T_2310 & _T_8 | ~_T_8 & _T_3867 : _T_3867;	// sequencer-master.scala:132:52, :184:52
      wire _T_3892 = io_op_bits_active_vfma ? _T_2311 & _T_8 | ~_T_8 & _T_3868 : _T_3868;	// sequencer-master.scala:132:52, :184:52
      wire _T_3893 = io_op_bits_active_vfma ? _T_2312 & _T_8 | ~_T_8 & _T_3869 : _T_3869;	// sequencer-master.scala:132:52, :184:52
      wire _T_3894 = io_op_bits_active_vfma ? _T_2313 & _T_8 | ~_T_8 & _T_3870 : _T_3870;	// sequencer-master.scala:132:52, :184:52
      wire _T_3895 = io_op_bits_active_vfma ? _T_2314 & _T_8 | ~_T_8 & _T_3871 : _T_3871;	// sequencer-master.scala:132:52, :184:52
      wire _T_3896 = io_op_bits_active_vfma ? _T_2315 & _T_8 | ~_T_8 & _T_3872 : _T_3872;	// sequencer-master.scala:132:52, :184:52
      wire _T_3897 = io_op_bits_active_vfma ? _T_2299 & _T_8 | ~_T_8 & _T_3873 : _T_3873;	// sequencer-master.scala:133:52, :185:52
      wire _T_3898 = io_op_bits_active_vfma ? _T_2300 & _T_8 | ~_T_8 & _T_3874 : _T_3874;	// sequencer-master.scala:133:52, :185:52
      wire _T_3899 = io_op_bits_active_vfma ? _T_2301 & _T_8 | ~_T_8 & _T_3875 : _T_3875;	// sequencer-master.scala:133:52, :185:52
      wire _T_3900 = io_op_bits_active_vfma ? _T_2302 & _T_8 | ~_T_8 & _T_3876 : _T_3876;	// sequencer-master.scala:133:52, :185:52
      wire _T_3901 = io_op_bits_active_vfma ? _T_2303 & _T_8 | ~_T_8 & _T_3877 : _T_3877;	// sequencer-master.scala:133:52, :185:52
      wire _T_3902 = io_op_bits_active_vfma ? _T_2304 & _T_8 | ~_T_8 & _T_3878 : _T_3878;	// sequencer-master.scala:133:52, :185:52
      wire _T_3903 = io_op_bits_active_vfma ? _T_2305 & _T_8 | ~_T_8 & _T_3879 : _T_3879;	// sequencer-master.scala:133:52, :185:52
      wire _T_3904 = io_op_bits_active_vfma ? _T_2306 & _T_8 | ~_T_8 & _T_3880 : _T_3880;	// sequencer-master.scala:133:52, :185:52
      wire _T_3905 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8 |
                ~_T_8 & _T_3881) : _T_3881;	// sequencer-master.scala:131:52, :183:52
      wire _T_3906 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8 |
                ~_T_8 & _T_3882) : _T_3882;	// sequencer-master.scala:131:52, :183:52
      wire _T_3907 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8 |
                ~_T_8 & _T_3883) : _T_3883;	// sequencer-master.scala:131:52, :183:52
      wire _T_3908 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8 |
                ~_T_8 & _T_3884) : _T_3884;	// sequencer-master.scala:131:52, :183:52
      wire _T_3909 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8 |
                ~_T_8 & _T_3885) : _T_3885;	// sequencer-master.scala:131:52, :183:52
      wire _T_3910 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8 |
                ~_T_8 & _T_3886) : _T_3886;	// sequencer-master.scala:131:52, :183:52
      wire _T_3911 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8 |
                ~_T_8 & _T_3887) : _T_3887;	// sequencer-master.scala:131:52, :183:52
      wire _T_3912 = io_op_bits_active_vfdiv ? ~_T_136 & (_T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8 |
                ~_T_8 & _T_3888) : _T_3888;	// sequencer-master.scala:131:52, :183:52
      wire _T_3913 = io_op_bits_active_vfdiv ? _T_2308 & _T_136 | ~_T_136 & (_T_2308 & _T_8 | ~_T_8 & _T_3889) :
                _T_3889;	// sequencer-master.scala:132:52, :184:52
      wire _T_3914 = io_op_bits_active_vfdiv ? _T_2309 & _T_136 | ~_T_136 & (_T_2309 & _T_8 | ~_T_8 & _T_3890) :
                _T_3890;	// sequencer-master.scala:132:52, :184:52
      wire _T_3915 = io_op_bits_active_vfdiv ? _T_2310 & _T_136 | ~_T_136 & (_T_2310 & _T_8 | ~_T_8 & _T_3891) :
                _T_3891;	// sequencer-master.scala:132:52, :184:52
      wire _T_3916 = io_op_bits_active_vfdiv ? _T_2311 & _T_136 | ~_T_136 & (_T_2311 & _T_8 | ~_T_8 & _T_3892) :
                _T_3892;	// sequencer-master.scala:132:52, :184:52
      wire _T_3917 = io_op_bits_active_vfdiv ? _T_2312 & _T_136 | ~_T_136 & (_T_2312 & _T_8 | ~_T_8 & _T_3893) :
                _T_3893;	// sequencer-master.scala:132:52, :184:52
      wire _T_3918 = io_op_bits_active_vfdiv ? _T_2313 & _T_136 | ~_T_136 & (_T_2313 & _T_8 | ~_T_8 & _T_3894) :
                _T_3894;	// sequencer-master.scala:132:52, :184:52
      wire _T_3919 = io_op_bits_active_vfdiv ? _T_2314 & _T_136 | ~_T_136 & (_T_2314 & _T_8 | ~_T_8 & _T_3895) :
                _T_3895;	// sequencer-master.scala:132:52, :184:52
      wire _T_3920 = io_op_bits_active_vfdiv ? _T_2315 & _T_136 | ~_T_136 & (_T_2315 & _T_8 | ~_T_8 & _T_3896) :
                _T_3896;	// sequencer-master.scala:132:52, :184:52
      wire _T_3921 = io_op_bits_active_vfdiv ? _T_2299 & _T_136 | ~_T_136 & (_T_2299 & _T_8 | ~_T_8 & _T_3897) :
                _T_3897;	// sequencer-master.scala:133:52, :185:52
      wire _T_3922 = io_op_bits_active_vfdiv ? _T_2300 & _T_136 | ~_T_136 & (_T_2300 & _T_8 | ~_T_8 & _T_3898) :
                _T_3898;	// sequencer-master.scala:133:52, :185:52
      wire _T_3923 = io_op_bits_active_vfdiv ? _T_2301 & _T_136 | ~_T_136 & (_T_2301 & _T_8 | ~_T_8 & _T_3899) :
                _T_3899;	// sequencer-master.scala:133:52, :185:52
      wire _T_3924 = io_op_bits_active_vfdiv ? _T_2302 & _T_136 | ~_T_136 & (_T_2302 & _T_8 | ~_T_8 & _T_3900) :
                _T_3900;	// sequencer-master.scala:133:52, :185:52
      wire _T_3925 = io_op_bits_active_vfdiv ? _T_2303 & _T_136 | ~_T_136 & (_T_2303 & _T_8 | ~_T_8 & _T_3901) :
                _T_3901;	// sequencer-master.scala:133:52, :185:52
      wire _T_3926 = io_op_bits_active_vfdiv ? _T_2304 & _T_136 | ~_T_136 & (_T_2304 & _T_8 | ~_T_8 & _T_3902) :
                _T_3902;	// sequencer-master.scala:133:52, :185:52
      wire _T_3927 = io_op_bits_active_vfdiv ? _T_2305 & _T_136 | ~_T_136 & (_T_2305 & _T_8 | ~_T_8 & _T_3903) :
                _T_3903;	// sequencer-master.scala:133:52, :185:52
      wire _T_3928 = io_op_bits_active_vfdiv ? _T_2306 & _T_136 | ~_T_136 & (_T_2306 & _T_8 | ~_T_8 & _T_3904) :
                _T_3904;	// sequencer-master.scala:133:52, :185:52
      wire _T_3929 = io_op_bits_active_vfcmp ? _T_2279 & _T_8 | _T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 &
                _T_3905 : _T_3905;	// sequencer-master.scala:131:52, :183:52
      wire _T_3930 = io_op_bits_active_vfcmp ? _T_2280 & _T_8 | _T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 &
                _T_3906 : _T_3906;	// sequencer-master.scala:131:52, :183:52
      wire _T_3931 = io_op_bits_active_vfcmp ? _T_2281 & _T_8 | _T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 &
                _T_3907 : _T_3907;	// sequencer-master.scala:131:52, :183:52
      wire _T_3932 = io_op_bits_active_vfcmp ? _T_2282 & _T_8 | _T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 &
                _T_3908 : _T_3908;	// sequencer-master.scala:131:52, :183:52
      wire _T_3933 = io_op_bits_active_vfcmp ? _T_2283 & _T_8 | _T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 &
                _T_3909 : _T_3909;	// sequencer-master.scala:131:52, :183:52
      wire _T_3934 = io_op_bits_active_vfcmp ? _T_2284 & _T_8 | _T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 &
                _T_3910 : _T_3910;	// sequencer-master.scala:131:52, :183:52
      wire _T_3935 = io_op_bits_active_vfcmp ? _T_2285 & _T_8 | _T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 &
                _T_3911 : _T_3911;	// sequencer-master.scala:131:52, :183:52
      wire _T_3936 = io_op_bits_active_vfcmp ? _T_2286 & _T_8 | _T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 &
                _T_3912 : _T_3912;	// sequencer-master.scala:131:52, :183:52
      wire _T_3937 = io_op_bits_active_vfcmp ? _T_2308 & _T_8 | ~_T_8 & _T_3913 : _T_3913;	// sequencer-master.scala:132:52, :184:52
      wire _T_3938 = io_op_bits_active_vfcmp ? _T_2309 & _T_8 | ~_T_8 & _T_3914 : _T_3914;	// sequencer-master.scala:132:52, :184:52
      wire _T_3939 = io_op_bits_active_vfcmp ? _T_2310 & _T_8 | ~_T_8 & _T_3915 : _T_3915;	// sequencer-master.scala:132:52, :184:52
      wire _T_3940 = io_op_bits_active_vfcmp ? _T_2311 & _T_8 | ~_T_8 & _T_3916 : _T_3916;	// sequencer-master.scala:132:52, :184:52
      wire _T_3941 = io_op_bits_active_vfcmp ? _T_2312 & _T_8 | ~_T_8 & _T_3917 : _T_3917;	// sequencer-master.scala:132:52, :184:52
      wire _T_3942 = io_op_bits_active_vfcmp ? _T_2313 & _T_8 | ~_T_8 & _T_3918 : _T_3918;	// sequencer-master.scala:132:52, :184:52
      wire _T_3943 = io_op_bits_active_vfcmp ? _T_2314 & _T_8 | ~_T_8 & _T_3919 : _T_3919;	// sequencer-master.scala:132:52, :184:52
      wire _T_3944 = io_op_bits_active_vfcmp ? _T_2315 & _T_8 | ~_T_8 & _T_3920 : _T_3920;	// sequencer-master.scala:132:52, :184:52
      wire _T_3945 = io_op_bits_active_vfcmp ? _T_2299 & _T_8 | ~_T_8 & _T_3921 : _T_3921;	// sequencer-master.scala:133:52, :185:52
      wire _T_3946 = io_op_bits_active_vfcmp ? _T_2300 & _T_8 | ~_T_8 & _T_3922 : _T_3922;	// sequencer-master.scala:133:52, :185:52
      wire _T_3947 = io_op_bits_active_vfcmp ? _T_2301 & _T_8 | ~_T_8 & _T_3923 : _T_3923;	// sequencer-master.scala:133:52, :185:52
      wire _T_3948 = io_op_bits_active_vfcmp ? _T_2302 & _T_8 | ~_T_8 & _T_3924 : _T_3924;	// sequencer-master.scala:133:52, :185:52
      wire _T_3949 = io_op_bits_active_vfcmp ? _T_2303 & _T_8 | ~_T_8 & _T_3925 : _T_3925;	// sequencer-master.scala:133:52, :185:52
      wire _T_3950 = io_op_bits_active_vfcmp ? _T_2304 & _T_8 | ~_T_8 & _T_3926 : _T_3926;	// sequencer-master.scala:133:52, :185:52
      wire _T_3951 = io_op_bits_active_vfcmp ? _T_2305 & _T_8 | ~_T_8 & _T_3927 : _T_3927;	// sequencer-master.scala:133:52, :185:52
      wire _T_3952 = io_op_bits_active_vfcmp ? _T_2306 & _T_8 | ~_T_8 & _T_3928 : _T_3928;	// sequencer-master.scala:133:52, :185:52
      wire _T_3953 = io_op_bits_active_vfconv ? _T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 & _T_3929 : _T_3929;	// sequencer-master.scala:131:52, :183:52
      wire _T_3954 = io_op_bits_active_vfconv ? _T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 & _T_3930 : _T_3930;	// sequencer-master.scala:131:52, :183:52
      wire _T_3955 = io_op_bits_active_vfconv ? _T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 & _T_3931 : _T_3931;	// sequencer-master.scala:131:52, :183:52
      wire _T_3956 = io_op_bits_active_vfconv ? _T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 & _T_3932 : _T_3932;	// sequencer-master.scala:131:52, :183:52
      wire _T_3957 = io_op_bits_active_vfconv ? _T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 & _T_3933 : _T_3933;	// sequencer-master.scala:131:52, :183:52
      wire _T_3958 = io_op_bits_active_vfconv ? _T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 & _T_3934 : _T_3934;	// sequencer-master.scala:131:52, :183:52
      wire _T_3959 = io_op_bits_active_vfconv ? _T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 & _T_3935 : _T_3935;	// sequencer-master.scala:131:52, :183:52
      wire _T_3960 = io_op_bits_active_vfconv ? _T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 & _T_3936 : _T_3936;	// sequencer-master.scala:131:52, :183:52
      wire _T_3961 = io_op_bits_active_vrpred ? _T_2238 & _T_8 | ~_T_8 & _T_3953 : _T_3953;	// sequencer-master.scala:131:52, :183:52
      wire _T_3962 = io_op_bits_active_vrpred ? _T_2242 & _T_8 | ~_T_8 & _T_3954 : _T_3954;	// sequencer-master.scala:131:52, :183:52
      wire _T_3963 = io_op_bits_active_vrpred ? _T_2246 & _T_8 | ~_T_8 & _T_3955 : _T_3955;	// sequencer-master.scala:131:52, :183:52
      wire _T_3964 = io_op_bits_active_vrpred ? _T_2250 & _T_8 | ~_T_8 & _T_3956 : _T_3956;	// sequencer-master.scala:131:52, :183:52
      wire _T_3965 = io_op_bits_active_vrpred ? _T_2254 & _T_8 | ~_T_8 & _T_3957 : _T_3957;	// sequencer-master.scala:131:52, :183:52
      wire _T_3966 = io_op_bits_active_vrpred ? _T_2258 & _T_8 | ~_T_8 & _T_3958 : _T_3958;	// sequencer-master.scala:131:52, :183:52
      wire _T_3967 = io_op_bits_active_vrpred ? _T_2262 & _T_8 | ~_T_8 & _T_3959 : _T_3959;	// sequencer-master.scala:131:52, :183:52
      wire _T_3968 = io_op_bits_active_vrpred ? _T_2266 & _T_8 | ~_T_8 & _T_3960 : _T_3960;	// sequencer-master.scala:131:52, :183:52
      wire _T_3969 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_8 | ~_T_8 & _T_3937 : _T_3937);	// sequencer-master.scala:132:52, :184:52
      wire _T_3970 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_8 | ~_T_8 & _T_3945 : _T_3945);	// sequencer-master.scala:133:52, :185:52
      wire _T_3971 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_8 | ~_T_8 & _T_3938 : _T_3938);	// sequencer-master.scala:132:52, :184:52
      wire _T_3972 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_8 | ~_T_8 & _T_3946 : _T_3946);	// sequencer-master.scala:133:52, :185:52
      wire _T_3973 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_8 | ~_T_8 & _T_3939 : _T_3939);	// sequencer-master.scala:132:52, :184:52
      wire _T_3974 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_8 | ~_T_8 & _T_3947 : _T_3947);	// sequencer-master.scala:133:52, :185:52
      wire _T_3975 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_8 | ~_T_8 & _T_3940 : _T_3940);	// sequencer-master.scala:132:52, :184:52
      wire _T_3976 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_8 | ~_T_8 & _T_3948 : _T_3948);	// sequencer-master.scala:133:52, :185:52
      wire _T_3977 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_8 | ~_T_8 & _T_3941 : _T_3941);	// sequencer-master.scala:132:52, :184:52
      wire _T_3978 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_8 | ~_T_8 & _T_3949 : _T_3949);	// sequencer-master.scala:133:52, :185:52
      wire _T_3979 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_8 | ~_T_8 & _T_3942 : _T_3942);	// sequencer-master.scala:132:52, :184:52
      wire _T_3980 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_8 | ~_T_8 & _T_3950 : _T_3950);	// sequencer-master.scala:133:52, :185:52
      wire _T_3981 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_8 | ~_T_8 & _T_3943 : _T_3943);	// sequencer-master.scala:132:52, :184:52
      wire _T_3982 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_8 | ~_T_8 & _T_3951 : _T_3951);	// sequencer-master.scala:133:52, :185:52
      wire _T_3983 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_8 | ~_T_8 & _T_3944 : _T_3944);	// sequencer-master.scala:132:52, :184:52
      wire _T_3984 = (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_8 | ~_T_8 & _T_3952 : _T_3952);	// sequencer-master.scala:133:52, :185:52
      wire _T_3985 = io_op_bits_active_vrfirst ? _T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 & _T_3961 : _T_3961;	// sequencer-master.scala:131:52, :183:52
      wire _T_3986 = io_op_bits_active_vrfirst ? _T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 & _T_3962 : _T_3962;	// sequencer-master.scala:131:52, :183:52
      wire _T_3987 = io_op_bits_active_vrfirst ? _T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 & _T_3963 : _T_3963;	// sequencer-master.scala:131:52, :183:52
      wire _T_3988 = io_op_bits_active_vrfirst ? _T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 & _T_3964 : _T_3964;	// sequencer-master.scala:131:52, :183:52
      wire _T_3989 = io_op_bits_active_vrfirst ? _T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 & _T_3965 : _T_3965;	// sequencer-master.scala:131:52, :183:52
      wire _T_3990 = io_op_bits_active_vrfirst ? _T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 & _T_3966 : _T_3966;	// sequencer-master.scala:131:52, :183:52
      wire _T_3991 = io_op_bits_active_vrfirst ? _T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 & _T_3967 : _T_3967;	// sequencer-master.scala:131:52, :183:52
      wire _T_3992 = io_op_bits_active_vrfirst ? _T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 & _T_3968 : _T_3968;	// sequencer-master.scala:131:52, :183:52
      wire _T_3993 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_132 | _T_2279 & _T_295 | _T_2238 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2269 & _T_8 | _T_2238 & _T_8 | ~_T_8 & _T_3985)) : _T_3985;	// sequencer-master.scala:131:52, :183:52
      wire _T_3994 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_133 | _T_2280 & _T_295 | _T_2242 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2270 & _T_8 | _T_2242 & _T_8 | ~_T_8 & _T_3986)) : _T_3986;	// sequencer-master.scala:131:52, :183:52
      wire _T_3995 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_134 | _T_2281 & _T_295 | _T_2246 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2271 & _T_8 | _T_2246 & _T_8 | ~_T_8 & _T_3987)) : _T_3987;	// sequencer-master.scala:131:52, :183:52
      wire _T_3996 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_135 | _T_2282 & _T_295 | _T_2250 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2272 & _T_8 | _T_2250 & _T_8 | ~_T_8 & _T_3988)) : _T_3988;	// sequencer-master.scala:131:52, :183:52
      wire _T_3997 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_136 | _T_2283 & _T_295 | _T_2254 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2273 & _T_8 | _T_2254 & _T_8 | ~_T_8 & _T_3989)) : _T_3989;	// sequencer-master.scala:131:52, :183:52
      wire _T_3998 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_137 | _T_2284 & _T_295 | _T_2258 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2274 & _T_8 | _T_2258 & _T_8 | ~_T_8 & _T_3990)) : _T_3990;	// sequencer-master.scala:131:52, :183:52
      wire _T_3999 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & _T_138 | _T_2285 & _T_295 | _T_2262 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2275 & _T_8 | _T_2262 & _T_8 | ~_T_8 & _T_3991)) : _T_3991;	// sequencer-master.scala:131:52, :183:52
      wire _T_4000 = io_op_bits_active_vamo ? ~_T_318 & (_T_295 & &_T_0 | _T_2286 & _T_295 | _T_2266 & _T_295 |
                ~_T_295 & ~_T_136 & (_T_2276 & _T_8 | _T_2266 & _T_8 | ~_T_8 & _T_3992)) : _T_3992;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4001 = io_op_bits_active_vamo ? _T_2308 & _T_318 | ~_T_318 & ~_T_295 & (_T_2308 & _T_136 | ~_T_136
                & ~_T_8 & _T_3969) : _T_3969;	// sequencer-master.scala:132:52, :184:52
      wire _T_4002 = io_op_bits_active_vamo ? _T_2309 & _T_318 | ~_T_318 & ~_T_295 & (_T_2309 & _T_136 | ~_T_136
                & ~_T_8 & _T_3971) : _T_3971;	// sequencer-master.scala:132:52, :184:52
      wire _T_4003 = io_op_bits_active_vamo ? _T_2310 & _T_318 | ~_T_318 & ~_T_295 & (_T_2310 & _T_136 | ~_T_136
                & ~_T_8 & _T_3973) : _T_3973;	// sequencer-master.scala:132:52, :184:52
      wire _T_4004 = io_op_bits_active_vamo ? _T_2311 & _T_318 | ~_T_318 & ~_T_295 & (_T_2311 & _T_136 | ~_T_136
                & ~_T_8 & _T_3975) : _T_3975;	// sequencer-master.scala:132:52, :184:52
      wire _T_4005 = io_op_bits_active_vamo ? _T_2312 & _T_318 | ~_T_318 & ~_T_295 & (_T_2312 & _T_136 | ~_T_136
                & ~_T_8 & _T_3977) : _T_3977;	// sequencer-master.scala:132:52, :184:52
      wire _T_4006 = io_op_bits_active_vamo ? _T_2313 & _T_318 | ~_T_318 & ~_T_295 & (_T_2313 & _T_136 | ~_T_136
                & ~_T_8 & _T_3979) : _T_3979;	// sequencer-master.scala:132:52, :184:52
      wire _T_4007 = io_op_bits_active_vamo ? _T_2314 & _T_318 | ~_T_318 & ~_T_295 & (_T_2314 & _T_136 | ~_T_136
                & ~_T_8 & _T_3981) : _T_3981;	// sequencer-master.scala:132:52, :184:52
      wire _T_4008 = io_op_bits_active_vamo ? _T_2315 & _T_318 | ~_T_318 & ~_T_295 & (_T_2315 & _T_136 | ~_T_136
                & ~_T_8 & _T_3983) : _T_3983;	// sequencer-master.scala:132:52, :184:52
      wire _T_4009 = io_op_bits_active_vamo ? _T_2299 & _T_318 | ~_T_318 & ~_T_295 & (_T_2299 & _T_136 | ~_T_136
                & ~_T_8 & _T_3970) : _T_3970;	// sequencer-master.scala:133:52, :185:52
      wire _T_4010 = io_op_bits_active_vamo ? _T_2300 & _T_318 | ~_T_318 & ~_T_295 & (_T_2300 & _T_136 | ~_T_136
                & ~_T_8 & _T_3972) : _T_3972;	// sequencer-master.scala:133:52, :185:52
      wire _T_4011 = io_op_bits_active_vamo ? _T_2301 & _T_318 | ~_T_318 & ~_T_295 & (_T_2301 & _T_136 | ~_T_136
                & ~_T_8 & _T_3974) : _T_3974;	// sequencer-master.scala:133:52, :185:52
      wire _T_4012 = io_op_bits_active_vamo ? _T_2302 & _T_318 | ~_T_318 & ~_T_295 & (_T_2302 & _T_136 | ~_T_136
                & ~_T_8 & _T_3976) : _T_3976;	// sequencer-master.scala:133:52, :185:52
      wire _T_4013 = io_op_bits_active_vamo ? _T_2303 & _T_318 | ~_T_318 & ~_T_295 & (_T_2303 & _T_136 | ~_T_136
                & ~_T_8 & _T_3978) : _T_3978;	// sequencer-master.scala:133:52, :185:52
      wire _T_4014 = io_op_bits_active_vamo ? _T_2304 & _T_318 | ~_T_318 & ~_T_295 & (_T_2304 & _T_136 | ~_T_136
                & ~_T_8 & _T_3980) : _T_3980;	// sequencer-master.scala:133:52, :185:52
      wire _T_4015 = io_op_bits_active_vamo ? _T_2305 & _T_318 | ~_T_318 & ~_T_295 & (_T_2305 & _T_136 | ~_T_136
                & ~_T_8 & _T_3982) : _T_3982;	// sequencer-master.scala:133:52, :185:52
      wire _T_4016 = io_op_bits_active_vamo ? _T_2306 & _T_318 | ~_T_318 & ~_T_295 & (_T_2306 & _T_136 | ~_T_136
                & ~_T_8 & _T_3984) : _T_3984;	// sequencer-master.scala:133:52, :185:52
      wire _T_4017 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2279 & _T_8 | _T_2238 & _T_8 | ~_T_8 &
                _T_3993) : _T_3993;	// sequencer-master.scala:131:52, :183:52
      wire _T_4018 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2280 & _T_8 | _T_2242 & _T_8 | ~_T_8 &
                _T_3994) : _T_3994;	// sequencer-master.scala:131:52, :183:52
      wire _T_4019 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2281 & _T_8 | _T_2246 & _T_8 | ~_T_8 &
                _T_3995) : _T_3995;	// sequencer-master.scala:131:52, :183:52
      wire _T_4020 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2282 & _T_8 | _T_2250 & _T_8 | ~_T_8 &
                _T_3996) : _T_3996;	// sequencer-master.scala:131:52, :183:52
      wire _T_4021 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2283 & _T_8 | _T_2254 & _T_8 | ~_T_8 &
                _T_3997) : _T_3997;	// sequencer-master.scala:131:52, :183:52
      wire _T_4022 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2284 & _T_8 | _T_2258 & _T_8 | ~_T_8 &
                _T_3998) : _T_3998;	// sequencer-master.scala:131:52, :183:52
      wire _T_4023 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2285 & _T_8 | _T_2262 & _T_8 | ~_T_8 &
                _T_3999) : _T_3999;	// sequencer-master.scala:131:52, :183:52
      wire _T_4024 = io_op_bits_active_vldx ? ~_T_295 & ~_T_136 & (_T_2286 & _T_8 | _T_2266 & _T_8 | ~_T_8 &
                _T_4000) : _T_4000;	// sequencer-master.scala:131:52, :183:52
      wire _T_4025 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2308 &
                _T_295 | ~_T_295 & (_T_2308 & _T_136 | ~_T_136 & ~_T_8 & _T_4001) : _T_4001);	// sequencer-master.scala:132:52, :184:52
      wire _T_4026 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2299 &
                _T_295 | ~_T_295 & (_T_2299 & _T_136 | ~_T_136 & ~_T_8 & _T_4009) : _T_4009);	// sequencer-master.scala:133:52, :185:52
      wire _T_4027 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2309 &
                _T_295 | ~_T_295 & (_T_2309 & _T_136 | ~_T_136 & ~_T_8 & _T_4002) : _T_4002);	// sequencer-master.scala:132:52, :184:52
      wire _T_4028 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2300 &
                _T_295 | ~_T_295 & (_T_2300 & _T_136 | ~_T_136 & ~_T_8 & _T_4010) : _T_4010);	// sequencer-master.scala:133:52, :185:52
      wire _T_4029 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2310 &
                _T_295 | ~_T_295 & (_T_2310 & _T_136 | ~_T_136 & ~_T_8 & _T_4003) : _T_4003);	// sequencer-master.scala:132:52, :184:52
      wire _T_4030 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2301 &
                _T_295 | ~_T_295 & (_T_2301 & _T_136 | ~_T_136 & ~_T_8 & _T_4011) : _T_4011);	// sequencer-master.scala:133:52, :185:52
      wire _T_4031 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2311 &
                _T_295 | ~_T_295 & (_T_2311 & _T_136 | ~_T_136 & ~_T_8 & _T_4004) : _T_4004);	// sequencer-master.scala:132:52, :184:52
      wire _T_4032 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2302 &
                _T_295 | ~_T_295 & (_T_2302 & _T_136 | ~_T_136 & ~_T_8 & _T_4012) : _T_4012);	// sequencer-master.scala:133:52, :185:52
      wire _T_4033 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2312 &
                _T_295 | ~_T_295 & (_T_2312 & _T_136 | ~_T_136 & ~_T_8 & _T_4005) : _T_4005);	// sequencer-master.scala:132:52, :184:52
      wire _T_4034 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2303 &
                _T_295 | ~_T_295 & (_T_2303 & _T_136 | ~_T_136 & ~_T_8 & _T_4013) : _T_4013);	// sequencer-master.scala:133:52, :185:52
      wire _T_4035 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2313 &
                _T_295 | ~_T_295 & (_T_2313 & _T_136 | ~_T_136 & ~_T_8 & _T_4006) : _T_4006);	// sequencer-master.scala:132:52, :184:52
      wire _T_4036 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2304 &
                _T_295 | ~_T_295 & (_T_2304 & _T_136 | ~_T_136 & ~_T_8 & _T_4014) : _T_4014);	// sequencer-master.scala:133:52, :185:52
      wire _T_4037 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2314 &
                _T_295 | ~_T_295 & (_T_2314 & _T_136 | ~_T_136 & ~_T_8 & _T_4007) : _T_4007);	// sequencer-master.scala:132:52, :184:52
      wire _T_4038 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2305 &
                _T_295 | ~_T_295 & (_T_2305 & _T_136 | ~_T_136 & ~_T_8 & _T_4015) : _T_4015);	// sequencer-master.scala:133:52, :185:52
      wire _T_4039 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2315 &
                _T_295 | ~_T_295 & (_T_2315 & _T_136 | ~_T_136 & ~_T_8 & _T_4008) : _T_4008);	// sequencer-master.scala:132:52, :184:52
      wire _T_4040 = (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vldx ? _T_2306 &
                _T_295 | ~_T_295 & (_T_2306 & _T_136 | ~_T_136 & ~_T_8 & _T_4016) : _T_4016);	// sequencer-master.scala:133:52, :185:52
      wire _T_4041 = io_op_bits_active_vstx ? _T_295 & _T_132 | _T_2299 & _T_295 | _T_2238 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2279 & _T_8 | _T_2238 & _T_8 | ~_T_8 & _T_4017) : _T_4017;	// sequencer-master.scala:131:52, :183:52
      wire _T_4042 = io_op_bits_active_vstx ? _T_295 & _T_133 | _T_2300 & _T_295 | _T_2242 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2280 & _T_8 | _T_2242 & _T_8 | ~_T_8 & _T_4018) : _T_4018;	// sequencer-master.scala:131:52, :183:52
      wire _T_4043 = io_op_bits_active_vstx ? _T_295 & _T_134 | _T_2301 & _T_295 | _T_2246 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2281 & _T_8 | _T_2246 & _T_8 | ~_T_8 & _T_4019) : _T_4019;	// sequencer-master.scala:131:52, :183:52
      wire _T_4044 = io_op_bits_active_vstx ? _T_295 & _T_135 | _T_2302 & _T_295 | _T_2250 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2282 & _T_8 | _T_2250 & _T_8 | ~_T_8 & _T_4020) : _T_4020;	// sequencer-master.scala:131:52, :183:52
      wire _T_4045 = io_op_bits_active_vstx ? _T_295 & _T_136 | _T_2303 & _T_295 | _T_2254 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2283 & _T_8 | _T_2254 & _T_8 | ~_T_8 & _T_4021) : _T_4021;	// sequencer-master.scala:131:52, :183:52
      wire _T_4046 = io_op_bits_active_vstx ? _T_295 & _T_137 | _T_2304 & _T_295 | _T_2258 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2284 & _T_8 | _T_2258 & _T_8 | ~_T_8 & _T_4022) : _T_4022;	// sequencer-master.scala:131:52, :183:52
      wire _T_4047 = io_op_bits_active_vstx ? _T_295 & _T_138 | _T_2305 & _T_295 | _T_2262 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2285 & _T_8 | _T_2262 & _T_8 | ~_T_8 & _T_4023) : _T_4023;	// sequencer-master.scala:131:52, :183:52
      wire _T_4048 = io_op_bits_active_vstx ? _T_295 & &_T_0 | _T_2306 & _T_295 | _T_2266 & _T_295 | ~_T_295 &
                ~_T_136 & (_T_2286 & _T_8 | _T_2266 & _T_8 | ~_T_8 & _T_4024) : _T_4024;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4049 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2238 & _T_8 | ~_T_8 & _T_4041) : _T_4041;	// sequencer-master.scala:131:52, :183:52
      wire _T_4050 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2242 & _T_8 | ~_T_8 & _T_4042) : _T_4042;	// sequencer-master.scala:131:52, :183:52
      wire _T_4051 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2246 & _T_8 | ~_T_8 & _T_4043) : _T_4043;	// sequencer-master.scala:131:52, :183:52
      wire _T_4052 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2250 & _T_8 | ~_T_8 & _T_4044) : _T_4044;	// sequencer-master.scala:131:52, :183:52
      wire _T_4053 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2254 & _T_8 | ~_T_8 & _T_4045) : _T_4045;	// sequencer-master.scala:131:52, :183:52
      wire _T_4054 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2258 & _T_8 | ~_T_8 & _T_4046) : _T_4046;	// sequencer-master.scala:131:52, :183:52
      wire _T_4055 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2262 & _T_8 | ~_T_8 & _T_4047) : _T_4047;	// sequencer-master.scala:131:52, :183:52
      wire _T_4056 = io_op_bits_active_vld ? ~_T_295 & ~_T_136 & (_T_2266 & _T_8 | ~_T_8 & _T_4048) : _T_4048;	// sequencer-master.scala:131:52, :183:52
      wire _T_4057 = io_op_bits_active_vint ? _T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 &
                e_5_raw_0 : e_5_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_4058 = io_op_bits_active_vint ? _T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 &
                e_5_raw_1 : e_5_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_4059 = io_op_bits_active_vint ? _T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 &
                e_5_raw_2 : e_5_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_4060 = io_op_bits_active_vint ? _T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 &
                e_5_raw_3 : e_5_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_4061 = io_op_bits_active_vint ? _T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 &
                e_5_raw_4 : e_5_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_4062 = io_op_bits_active_vint ? _T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 &
                e_5_raw_5 : e_5_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_4063 = io_op_bits_active_vint ? _T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 &
                e_5_raw_6 : e_5_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_4064 = io_op_bits_active_vint ? _T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 &
                e_5_raw_7 : e_5_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_4065 = io_op_bits_active_vint ? _T_2308 & _T_9 | ~_T_9 & e_5_war_0 : e_5_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_4066 = io_op_bits_active_vint ? _T_2309 & _T_9 | ~_T_9 & e_5_war_1 : e_5_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_4067 = io_op_bits_active_vint ? _T_2310 & _T_9 | ~_T_9 & e_5_war_2 : e_5_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_4068 = io_op_bits_active_vint ? _T_2311 & _T_9 | ~_T_9 & e_5_war_3 : e_5_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_4069 = io_op_bits_active_vint ? _T_2312 & _T_9 | ~_T_9 & e_5_war_4 : e_5_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_4070 = io_op_bits_active_vint ? _T_2313 & _T_9 | ~_T_9 & e_5_war_5 : e_5_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_4071 = io_op_bits_active_vint ? _T_2314 & _T_9 | ~_T_9 & e_5_war_6 : e_5_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_4072 = io_op_bits_active_vint ? _T_2315 & _T_9 | ~_T_9 & e_5_war_7 : e_5_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_4073 = io_op_bits_active_vint ? _T_2299 & _T_9 | ~_T_9 & e_5_waw_0 : e_5_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_4074 = io_op_bits_active_vint ? _T_2300 & _T_9 | ~_T_9 & e_5_waw_1 : e_5_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_4075 = io_op_bits_active_vint ? _T_2301 & _T_9 | ~_T_9 & e_5_waw_2 : e_5_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_4076 = io_op_bits_active_vint ? _T_2302 & _T_9 | ~_T_9 & e_5_waw_3 : e_5_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_4077 = io_op_bits_active_vint ? _T_2303 & _T_9 | ~_T_9 & e_5_waw_4 : e_5_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_4078 = io_op_bits_active_vint ? _T_2304 & _T_9 | ~_T_9 & e_5_waw_5 : e_5_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_4079 = io_op_bits_active_vint ? _T_2305 & _T_9 | ~_T_9 & e_5_waw_6 : e_5_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_4080 = io_op_bits_active_vint ? _T_2306 & _T_9 | ~_T_9 & e_5_waw_7 : e_5_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_4081 = io_op_bits_active_vipred ? _T_2289 & _T_9 | _T_2279 & _T_9 | _T_2269 & _T_9 | ~_T_9 &
                _T_4057 : _T_4057;	// sequencer-master.scala:131:52, :183:52
      wire _T_4082 = io_op_bits_active_vipred ? _T_2290 & _T_9 | _T_2280 & _T_9 | _T_2270 & _T_9 | ~_T_9 &
                _T_4058 : _T_4058;	// sequencer-master.scala:131:52, :183:52
      wire _T_4083 = io_op_bits_active_vipred ? _T_2291 & _T_9 | _T_2281 & _T_9 | _T_2271 & _T_9 | ~_T_9 &
                _T_4059 : _T_4059;	// sequencer-master.scala:131:52, :183:52
      wire _T_4084 = io_op_bits_active_vipred ? _T_2292 & _T_9 | _T_2282 & _T_9 | _T_2272 & _T_9 | ~_T_9 &
                _T_4060 : _T_4060;	// sequencer-master.scala:131:52, :183:52
      wire _T_4085 = io_op_bits_active_vipred ? _T_2293 & _T_9 | _T_2283 & _T_9 | _T_2273 & _T_9 | ~_T_9 &
                _T_4061 : _T_4061;	// sequencer-master.scala:131:52, :183:52
      wire _T_4086 = io_op_bits_active_vipred ? _T_2294 & _T_9 | _T_2284 & _T_9 | _T_2274 & _T_9 | ~_T_9 &
                _T_4062 : _T_4062;	// sequencer-master.scala:131:52, :183:52
      wire _T_4087 = io_op_bits_active_vipred ? _T_2295 & _T_9 | _T_2285 & _T_9 | _T_2275 & _T_9 | ~_T_9 &
                _T_4063 : _T_4063;	// sequencer-master.scala:131:52, :183:52
      wire _T_4088 = io_op_bits_active_vipred ? _T_2296 & _T_9 | _T_2286 & _T_9 | _T_2276 & _T_9 | ~_T_9 &
                _T_4064 : _T_4064;	// sequencer-master.scala:131:52, :183:52
      wire _T_4089 = io_op_bits_active_vipred ? _T_2308 & _T_9 | ~_T_9 & _T_4065 : _T_4065;	// sequencer-master.scala:132:52, :184:52
      wire _T_4090 = io_op_bits_active_vipred ? _T_2309 & _T_9 | ~_T_9 & _T_4066 : _T_4066;	// sequencer-master.scala:132:52, :184:52
      wire _T_4091 = io_op_bits_active_vipred ? _T_2310 & _T_9 | ~_T_9 & _T_4067 : _T_4067;	// sequencer-master.scala:132:52, :184:52
      wire _T_4092 = io_op_bits_active_vipred ? _T_2311 & _T_9 | ~_T_9 & _T_4068 : _T_4068;	// sequencer-master.scala:132:52, :184:52
      wire _T_4093 = io_op_bits_active_vipred ? _T_2312 & _T_9 | ~_T_9 & _T_4069 : _T_4069;	// sequencer-master.scala:132:52, :184:52
      wire _T_4094 = io_op_bits_active_vipred ? _T_2313 & _T_9 | ~_T_9 & _T_4070 : _T_4070;	// sequencer-master.scala:132:52, :184:52
      wire _T_4095 = io_op_bits_active_vipred ? _T_2314 & _T_9 | ~_T_9 & _T_4071 : _T_4071;	// sequencer-master.scala:132:52, :184:52
      wire _T_4096 = io_op_bits_active_vipred ? _T_2315 & _T_9 | ~_T_9 & _T_4072 : _T_4072;	// sequencer-master.scala:132:52, :184:52
      wire _T_4097 = io_op_bits_active_vipred ? _T_2299 & _T_9 | ~_T_9 & _T_4073 : _T_4073;	// sequencer-master.scala:133:52, :185:52
      wire _T_4098 = io_op_bits_active_vipred ? _T_2300 & _T_9 | ~_T_9 & _T_4074 : _T_4074;	// sequencer-master.scala:133:52, :185:52
      wire _T_4099 = io_op_bits_active_vipred ? _T_2301 & _T_9 | ~_T_9 & _T_4075 : _T_4075;	// sequencer-master.scala:133:52, :185:52
      wire _T_4100 = io_op_bits_active_vipred ? _T_2302 & _T_9 | ~_T_9 & _T_4076 : _T_4076;	// sequencer-master.scala:133:52, :185:52
      wire _T_4101 = io_op_bits_active_vipred ? _T_2303 & _T_9 | ~_T_9 & _T_4077 : _T_4077;	// sequencer-master.scala:133:52, :185:52
      wire _T_4102 = io_op_bits_active_vipred ? _T_2304 & _T_9 | ~_T_9 & _T_4078 : _T_4078;	// sequencer-master.scala:133:52, :185:52
      wire _T_4103 = io_op_bits_active_vipred ? _T_2305 & _T_9 | ~_T_9 & _T_4079 : _T_4079;	// sequencer-master.scala:133:52, :185:52
      wire _T_4104 = io_op_bits_active_vipred ? _T_2306 & _T_9 | ~_T_9 & _T_4080 : _T_4080;	// sequencer-master.scala:133:52, :185:52
      wire _T_4105 = io_op_bits_active_vimul ? _T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 &
                _T_4081 : _T_4081;	// sequencer-master.scala:131:52, :183:52
      wire _T_4106 = io_op_bits_active_vimul ? _T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 &
                _T_4082 : _T_4082;	// sequencer-master.scala:131:52, :183:52
      wire _T_4107 = io_op_bits_active_vimul ? _T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 &
                _T_4083 : _T_4083;	// sequencer-master.scala:131:52, :183:52
      wire _T_4108 = io_op_bits_active_vimul ? _T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 &
                _T_4084 : _T_4084;	// sequencer-master.scala:131:52, :183:52
      wire _T_4109 = io_op_bits_active_vimul ? _T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 &
                _T_4085 : _T_4085;	// sequencer-master.scala:131:52, :183:52
      wire _T_4110 = io_op_bits_active_vimul ? _T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 &
                _T_4086 : _T_4086;	// sequencer-master.scala:131:52, :183:52
      wire _T_4111 = io_op_bits_active_vimul ? _T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 &
                _T_4087 : _T_4087;	// sequencer-master.scala:131:52, :183:52
      wire _T_4112 = io_op_bits_active_vimul ? _T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 &
                _T_4088 : _T_4088;	// sequencer-master.scala:131:52, :183:52
      wire _T_4113 = io_op_bits_active_vimul ? _T_2308 & _T_9 | ~_T_9 & _T_4089 : _T_4089;	// sequencer-master.scala:132:52, :184:52
      wire _T_4114 = io_op_bits_active_vimul ? _T_2309 & _T_9 | ~_T_9 & _T_4090 : _T_4090;	// sequencer-master.scala:132:52, :184:52
      wire _T_4115 = io_op_bits_active_vimul ? _T_2310 & _T_9 | ~_T_9 & _T_4091 : _T_4091;	// sequencer-master.scala:132:52, :184:52
      wire _T_4116 = io_op_bits_active_vimul ? _T_2311 & _T_9 | ~_T_9 & _T_4092 : _T_4092;	// sequencer-master.scala:132:52, :184:52
      wire _T_4117 = io_op_bits_active_vimul ? _T_2312 & _T_9 | ~_T_9 & _T_4093 : _T_4093;	// sequencer-master.scala:132:52, :184:52
      wire _T_4118 = io_op_bits_active_vimul ? _T_2313 & _T_9 | ~_T_9 & _T_4094 : _T_4094;	// sequencer-master.scala:132:52, :184:52
      wire _T_4119 = io_op_bits_active_vimul ? _T_2314 & _T_9 | ~_T_9 & _T_4095 : _T_4095;	// sequencer-master.scala:132:52, :184:52
      wire _T_4120 = io_op_bits_active_vimul ? _T_2315 & _T_9 | ~_T_9 & _T_4096 : _T_4096;	// sequencer-master.scala:132:52, :184:52
      wire _T_4121 = io_op_bits_active_vimul ? _T_2299 & _T_9 | ~_T_9 & _T_4097 : _T_4097;	// sequencer-master.scala:133:52, :185:52
      wire _T_4122 = io_op_bits_active_vimul ? _T_2300 & _T_9 | ~_T_9 & _T_4098 : _T_4098;	// sequencer-master.scala:133:52, :185:52
      wire _T_4123 = io_op_bits_active_vimul ? _T_2301 & _T_9 | ~_T_9 & _T_4099 : _T_4099;	// sequencer-master.scala:133:52, :185:52
      wire _T_4124 = io_op_bits_active_vimul ? _T_2302 & _T_9 | ~_T_9 & _T_4100 : _T_4100;	// sequencer-master.scala:133:52, :185:52
      wire _T_4125 = io_op_bits_active_vimul ? _T_2303 & _T_9 | ~_T_9 & _T_4101 : _T_4101;	// sequencer-master.scala:133:52, :185:52
      wire _T_4126 = io_op_bits_active_vimul ? _T_2304 & _T_9 | ~_T_9 & _T_4102 : _T_4102;	// sequencer-master.scala:133:52, :185:52
      wire _T_4127 = io_op_bits_active_vimul ? _T_2305 & _T_9 | ~_T_9 & _T_4103 : _T_4103;	// sequencer-master.scala:133:52, :185:52
      wire _T_4128 = io_op_bits_active_vimul ? _T_2306 & _T_9 | ~_T_9 & _T_4104 : _T_4104;	// sequencer-master.scala:133:52, :185:52
      wire _T_4129 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9 |
                ~_T_9 & _T_4105) : _T_4105;	// sequencer-master.scala:131:52, :183:52
      wire _T_4130 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9 |
                ~_T_9 & _T_4106) : _T_4106;	// sequencer-master.scala:131:52, :183:52
      wire _T_4131 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9 |
                ~_T_9 & _T_4107) : _T_4107;	// sequencer-master.scala:131:52, :183:52
      wire _T_4132 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9 |
                ~_T_9 & _T_4108) : _T_4108;	// sequencer-master.scala:131:52, :183:52
      wire _T_4133 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9 |
                ~_T_9 & _T_4109) : _T_4109;	// sequencer-master.scala:131:52, :183:52
      wire _T_4134 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9 |
                ~_T_9 & _T_4110) : _T_4110;	// sequencer-master.scala:131:52, :183:52
      wire _T_4135 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9 |
                ~_T_9 & _T_4111) : _T_4111;	// sequencer-master.scala:131:52, :183:52
      wire _T_4136 = io_op_bits_active_vidiv ? ~_T_137 & (_T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9 |
                ~_T_9 & _T_4112) : _T_4112;	// sequencer-master.scala:131:52, :183:52
      wire _T_4137 = io_op_bits_active_vidiv ? _T_2308 & _T_137 | ~_T_137 & (_T_2308 & _T_9 | ~_T_9 & _T_4113) :
                _T_4113;	// sequencer-master.scala:132:52, :184:52
      wire _T_4138 = io_op_bits_active_vidiv ? _T_2309 & _T_137 | ~_T_137 & (_T_2309 & _T_9 | ~_T_9 & _T_4114) :
                _T_4114;	// sequencer-master.scala:132:52, :184:52
      wire _T_4139 = io_op_bits_active_vidiv ? _T_2310 & _T_137 | ~_T_137 & (_T_2310 & _T_9 | ~_T_9 & _T_4115) :
                _T_4115;	// sequencer-master.scala:132:52, :184:52
      wire _T_4140 = io_op_bits_active_vidiv ? _T_2311 & _T_137 | ~_T_137 & (_T_2311 & _T_9 | ~_T_9 & _T_4116) :
                _T_4116;	// sequencer-master.scala:132:52, :184:52
      wire _T_4141 = io_op_bits_active_vidiv ? _T_2312 & _T_137 | ~_T_137 & (_T_2312 & _T_9 | ~_T_9 & _T_4117) :
                _T_4117;	// sequencer-master.scala:132:52, :184:52
      wire _T_4142 = io_op_bits_active_vidiv ? _T_2313 & _T_137 | ~_T_137 & (_T_2313 & _T_9 | ~_T_9 & _T_4118) :
                _T_4118;	// sequencer-master.scala:132:52, :184:52
      wire _T_4143 = io_op_bits_active_vidiv ? _T_2314 & _T_137 | ~_T_137 & (_T_2314 & _T_9 | ~_T_9 & _T_4119) :
                _T_4119;	// sequencer-master.scala:132:52, :184:52
      wire _T_4144 = io_op_bits_active_vidiv ? _T_2315 & _T_137 | ~_T_137 & (_T_2315 & _T_9 | ~_T_9 & _T_4120) :
                _T_4120;	// sequencer-master.scala:132:52, :184:52
      wire _T_4145 = io_op_bits_active_vidiv ? _T_2299 & _T_137 | ~_T_137 & (_T_2299 & _T_9 | ~_T_9 & _T_4121) :
                _T_4121;	// sequencer-master.scala:133:52, :185:52
      wire _T_4146 = io_op_bits_active_vidiv ? _T_2300 & _T_137 | ~_T_137 & (_T_2300 & _T_9 | ~_T_9 & _T_4122) :
                _T_4122;	// sequencer-master.scala:133:52, :185:52
      wire _T_4147 = io_op_bits_active_vidiv ? _T_2301 & _T_137 | ~_T_137 & (_T_2301 & _T_9 | ~_T_9 & _T_4123) :
                _T_4123;	// sequencer-master.scala:133:52, :185:52
      wire _T_4148 = io_op_bits_active_vidiv ? _T_2302 & _T_137 | ~_T_137 & (_T_2302 & _T_9 | ~_T_9 & _T_4124) :
                _T_4124;	// sequencer-master.scala:133:52, :185:52
      wire _T_4149 = io_op_bits_active_vidiv ? _T_2303 & _T_137 | ~_T_137 & (_T_2303 & _T_9 | ~_T_9 & _T_4125) :
                _T_4125;	// sequencer-master.scala:133:52, :185:52
      wire _T_4150 = io_op_bits_active_vidiv ? _T_2304 & _T_137 | ~_T_137 & (_T_2304 & _T_9 | ~_T_9 & _T_4126) :
                _T_4126;	// sequencer-master.scala:133:52, :185:52
      wire _T_4151 = io_op_bits_active_vidiv ? _T_2305 & _T_137 | ~_T_137 & (_T_2305 & _T_9 | ~_T_9 & _T_4127) :
                _T_4127;	// sequencer-master.scala:133:52, :185:52
      wire _T_4152 = io_op_bits_active_vidiv ? _T_2306 & _T_137 | ~_T_137 & (_T_2306 & _T_9 | ~_T_9 & _T_4128) :
                _T_4128;	// sequencer-master.scala:133:52, :185:52
      wire _T_4153 = io_op_bits_active_vfma ? _T_2289 & _T_9 | _T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9
                | ~_T_9 & _T_4129 : _T_4129;	// sequencer-master.scala:131:52, :183:52
      wire _T_4154 = io_op_bits_active_vfma ? _T_2290 & _T_9 | _T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9
                | ~_T_9 & _T_4130 : _T_4130;	// sequencer-master.scala:131:52, :183:52
      wire _T_4155 = io_op_bits_active_vfma ? _T_2291 & _T_9 | _T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9
                | ~_T_9 & _T_4131 : _T_4131;	// sequencer-master.scala:131:52, :183:52
      wire _T_4156 = io_op_bits_active_vfma ? _T_2292 & _T_9 | _T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9
                | ~_T_9 & _T_4132 : _T_4132;	// sequencer-master.scala:131:52, :183:52
      wire _T_4157 = io_op_bits_active_vfma ? _T_2293 & _T_9 | _T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9
                | ~_T_9 & _T_4133 : _T_4133;	// sequencer-master.scala:131:52, :183:52
      wire _T_4158 = io_op_bits_active_vfma ? _T_2294 & _T_9 | _T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9
                | ~_T_9 & _T_4134 : _T_4134;	// sequencer-master.scala:131:52, :183:52
      wire _T_4159 = io_op_bits_active_vfma ? _T_2295 & _T_9 | _T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9
                | ~_T_9 & _T_4135 : _T_4135;	// sequencer-master.scala:131:52, :183:52
      wire _T_4160 = io_op_bits_active_vfma ? _T_2296 & _T_9 | _T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9
                | ~_T_9 & _T_4136 : _T_4136;	// sequencer-master.scala:131:52, :183:52
      wire _T_4161 = io_op_bits_active_vfma ? _T_2308 & _T_9 | ~_T_9 & _T_4137 : _T_4137;	// sequencer-master.scala:132:52, :184:52
      wire _T_4162 = io_op_bits_active_vfma ? _T_2309 & _T_9 | ~_T_9 & _T_4138 : _T_4138;	// sequencer-master.scala:132:52, :184:52
      wire _T_4163 = io_op_bits_active_vfma ? _T_2310 & _T_9 | ~_T_9 & _T_4139 : _T_4139;	// sequencer-master.scala:132:52, :184:52
      wire _T_4164 = io_op_bits_active_vfma ? _T_2311 & _T_9 | ~_T_9 & _T_4140 : _T_4140;	// sequencer-master.scala:132:52, :184:52
      wire _T_4165 = io_op_bits_active_vfma ? _T_2312 & _T_9 | ~_T_9 & _T_4141 : _T_4141;	// sequencer-master.scala:132:52, :184:52
      wire _T_4166 = io_op_bits_active_vfma ? _T_2313 & _T_9 | ~_T_9 & _T_4142 : _T_4142;	// sequencer-master.scala:132:52, :184:52
      wire _T_4167 = io_op_bits_active_vfma ? _T_2314 & _T_9 | ~_T_9 & _T_4143 : _T_4143;	// sequencer-master.scala:132:52, :184:52
      wire _T_4168 = io_op_bits_active_vfma ? _T_2315 & _T_9 | ~_T_9 & _T_4144 : _T_4144;	// sequencer-master.scala:132:52, :184:52
      wire _T_4169 = io_op_bits_active_vfma ? _T_2299 & _T_9 | ~_T_9 & _T_4145 : _T_4145;	// sequencer-master.scala:133:52, :185:52
      wire _T_4170 = io_op_bits_active_vfma ? _T_2300 & _T_9 | ~_T_9 & _T_4146 : _T_4146;	// sequencer-master.scala:133:52, :185:52
      wire _T_4171 = io_op_bits_active_vfma ? _T_2301 & _T_9 | ~_T_9 & _T_4147 : _T_4147;	// sequencer-master.scala:133:52, :185:52
      wire _T_4172 = io_op_bits_active_vfma ? _T_2302 & _T_9 | ~_T_9 & _T_4148 : _T_4148;	// sequencer-master.scala:133:52, :185:52
      wire _T_4173 = io_op_bits_active_vfma ? _T_2303 & _T_9 | ~_T_9 & _T_4149 : _T_4149;	// sequencer-master.scala:133:52, :185:52
      wire _T_4174 = io_op_bits_active_vfma ? _T_2304 & _T_9 | ~_T_9 & _T_4150 : _T_4150;	// sequencer-master.scala:133:52, :185:52
      wire _T_4175 = io_op_bits_active_vfma ? _T_2305 & _T_9 | ~_T_9 & _T_4151 : _T_4151;	// sequencer-master.scala:133:52, :185:52
      wire _T_4176 = io_op_bits_active_vfma ? _T_2306 & _T_9 | ~_T_9 & _T_4152 : _T_4152;	// sequencer-master.scala:133:52, :185:52
      wire _T_4177 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9 |
                ~_T_9 & _T_4153) : _T_4153;	// sequencer-master.scala:131:52, :183:52
      wire _T_4178 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9 |
                ~_T_9 & _T_4154) : _T_4154;	// sequencer-master.scala:131:52, :183:52
      wire _T_4179 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9 |
                ~_T_9 & _T_4155) : _T_4155;	// sequencer-master.scala:131:52, :183:52
      wire _T_4180 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9 |
                ~_T_9 & _T_4156) : _T_4156;	// sequencer-master.scala:131:52, :183:52
      wire _T_4181 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9 |
                ~_T_9 & _T_4157) : _T_4157;	// sequencer-master.scala:131:52, :183:52
      wire _T_4182 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9 |
                ~_T_9 & _T_4158) : _T_4158;	// sequencer-master.scala:131:52, :183:52
      wire _T_4183 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9 |
                ~_T_9 & _T_4159) : _T_4159;	// sequencer-master.scala:131:52, :183:52
      wire _T_4184 = io_op_bits_active_vfdiv ? ~_T_137 & (_T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9 |
                ~_T_9 & _T_4160) : _T_4160;	// sequencer-master.scala:131:52, :183:52
      wire _T_4185 = io_op_bits_active_vfdiv ? _T_2308 & _T_137 | ~_T_137 & (_T_2308 & _T_9 | ~_T_9 & _T_4161) :
                _T_4161;	// sequencer-master.scala:132:52, :184:52
      wire _T_4186 = io_op_bits_active_vfdiv ? _T_2309 & _T_137 | ~_T_137 & (_T_2309 & _T_9 | ~_T_9 & _T_4162) :
                _T_4162;	// sequencer-master.scala:132:52, :184:52
      wire _T_4187 = io_op_bits_active_vfdiv ? _T_2310 & _T_137 | ~_T_137 & (_T_2310 & _T_9 | ~_T_9 & _T_4163) :
                _T_4163;	// sequencer-master.scala:132:52, :184:52
      wire _T_4188 = io_op_bits_active_vfdiv ? _T_2311 & _T_137 | ~_T_137 & (_T_2311 & _T_9 | ~_T_9 & _T_4164) :
                _T_4164;	// sequencer-master.scala:132:52, :184:52
      wire _T_4189 = io_op_bits_active_vfdiv ? _T_2312 & _T_137 | ~_T_137 & (_T_2312 & _T_9 | ~_T_9 & _T_4165) :
                _T_4165;	// sequencer-master.scala:132:52, :184:52
      wire _T_4190 = io_op_bits_active_vfdiv ? _T_2313 & _T_137 | ~_T_137 & (_T_2313 & _T_9 | ~_T_9 & _T_4166) :
                _T_4166;	// sequencer-master.scala:132:52, :184:52
      wire _T_4191 = io_op_bits_active_vfdiv ? _T_2314 & _T_137 | ~_T_137 & (_T_2314 & _T_9 | ~_T_9 & _T_4167) :
                _T_4167;	// sequencer-master.scala:132:52, :184:52
      wire _T_4192 = io_op_bits_active_vfdiv ? _T_2315 & _T_137 | ~_T_137 & (_T_2315 & _T_9 | ~_T_9 & _T_4168) :
                _T_4168;	// sequencer-master.scala:132:52, :184:52
      wire _T_4193 = io_op_bits_active_vfdiv ? _T_2299 & _T_137 | ~_T_137 & (_T_2299 & _T_9 | ~_T_9 & _T_4169) :
                _T_4169;	// sequencer-master.scala:133:52, :185:52
      wire _T_4194 = io_op_bits_active_vfdiv ? _T_2300 & _T_137 | ~_T_137 & (_T_2300 & _T_9 | ~_T_9 & _T_4170) :
                _T_4170;	// sequencer-master.scala:133:52, :185:52
      wire _T_4195 = io_op_bits_active_vfdiv ? _T_2301 & _T_137 | ~_T_137 & (_T_2301 & _T_9 | ~_T_9 & _T_4171) :
                _T_4171;	// sequencer-master.scala:133:52, :185:52
      wire _T_4196 = io_op_bits_active_vfdiv ? _T_2302 & _T_137 | ~_T_137 & (_T_2302 & _T_9 | ~_T_9 & _T_4172) :
                _T_4172;	// sequencer-master.scala:133:52, :185:52
      wire _T_4197 = io_op_bits_active_vfdiv ? _T_2303 & _T_137 | ~_T_137 & (_T_2303 & _T_9 | ~_T_9 & _T_4173) :
                _T_4173;	// sequencer-master.scala:133:52, :185:52
      wire _T_4198 = io_op_bits_active_vfdiv ? _T_2304 & _T_137 | ~_T_137 & (_T_2304 & _T_9 | ~_T_9 & _T_4174) :
                _T_4174;	// sequencer-master.scala:133:52, :185:52
      wire _T_4199 = io_op_bits_active_vfdiv ? _T_2305 & _T_137 | ~_T_137 & (_T_2305 & _T_9 | ~_T_9 & _T_4175) :
                _T_4175;	// sequencer-master.scala:133:52, :185:52
      wire _T_4200 = io_op_bits_active_vfdiv ? _T_2306 & _T_137 | ~_T_137 & (_T_2306 & _T_9 | ~_T_9 & _T_4176) :
                _T_4176;	// sequencer-master.scala:133:52, :185:52
      wire _T_4201 = io_op_bits_active_vfcmp ? _T_2279 & _T_9 | _T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 &
                _T_4177 : _T_4177;	// sequencer-master.scala:131:52, :183:52
      wire _T_4202 = io_op_bits_active_vfcmp ? _T_2280 & _T_9 | _T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 &
                _T_4178 : _T_4178;	// sequencer-master.scala:131:52, :183:52
      wire _T_4203 = io_op_bits_active_vfcmp ? _T_2281 & _T_9 | _T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 &
                _T_4179 : _T_4179;	// sequencer-master.scala:131:52, :183:52
      wire _T_4204 = io_op_bits_active_vfcmp ? _T_2282 & _T_9 | _T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 &
                _T_4180 : _T_4180;	// sequencer-master.scala:131:52, :183:52
      wire _T_4205 = io_op_bits_active_vfcmp ? _T_2283 & _T_9 | _T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 &
                _T_4181 : _T_4181;	// sequencer-master.scala:131:52, :183:52
      wire _T_4206 = io_op_bits_active_vfcmp ? _T_2284 & _T_9 | _T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 &
                _T_4182 : _T_4182;	// sequencer-master.scala:131:52, :183:52
      wire _T_4207 = io_op_bits_active_vfcmp ? _T_2285 & _T_9 | _T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 &
                _T_4183 : _T_4183;	// sequencer-master.scala:131:52, :183:52
      wire _T_4208 = io_op_bits_active_vfcmp ? _T_2286 & _T_9 | _T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 &
                _T_4184 : _T_4184;	// sequencer-master.scala:131:52, :183:52
      wire _T_4209 = io_op_bits_active_vfcmp ? _T_2308 & _T_9 | ~_T_9 & _T_4185 : _T_4185;	// sequencer-master.scala:132:52, :184:52
      wire _T_4210 = io_op_bits_active_vfcmp ? _T_2309 & _T_9 | ~_T_9 & _T_4186 : _T_4186;	// sequencer-master.scala:132:52, :184:52
      wire _T_4211 = io_op_bits_active_vfcmp ? _T_2310 & _T_9 | ~_T_9 & _T_4187 : _T_4187;	// sequencer-master.scala:132:52, :184:52
      wire _T_4212 = io_op_bits_active_vfcmp ? _T_2311 & _T_9 | ~_T_9 & _T_4188 : _T_4188;	// sequencer-master.scala:132:52, :184:52
      wire _T_4213 = io_op_bits_active_vfcmp ? _T_2312 & _T_9 | ~_T_9 & _T_4189 : _T_4189;	// sequencer-master.scala:132:52, :184:52
      wire _T_4214 = io_op_bits_active_vfcmp ? _T_2313 & _T_9 | ~_T_9 & _T_4190 : _T_4190;	// sequencer-master.scala:132:52, :184:52
      wire _T_4215 = io_op_bits_active_vfcmp ? _T_2314 & _T_9 | ~_T_9 & _T_4191 : _T_4191;	// sequencer-master.scala:132:52, :184:52
      wire _T_4216 = io_op_bits_active_vfcmp ? _T_2315 & _T_9 | ~_T_9 & _T_4192 : _T_4192;	// sequencer-master.scala:132:52, :184:52
      wire _T_4217 = io_op_bits_active_vfcmp ? _T_2299 & _T_9 | ~_T_9 & _T_4193 : _T_4193;	// sequencer-master.scala:133:52, :185:52
      wire _T_4218 = io_op_bits_active_vfcmp ? _T_2300 & _T_9 | ~_T_9 & _T_4194 : _T_4194;	// sequencer-master.scala:133:52, :185:52
      wire _T_4219 = io_op_bits_active_vfcmp ? _T_2301 & _T_9 | ~_T_9 & _T_4195 : _T_4195;	// sequencer-master.scala:133:52, :185:52
      wire _T_4220 = io_op_bits_active_vfcmp ? _T_2302 & _T_9 | ~_T_9 & _T_4196 : _T_4196;	// sequencer-master.scala:133:52, :185:52
      wire _T_4221 = io_op_bits_active_vfcmp ? _T_2303 & _T_9 | ~_T_9 & _T_4197 : _T_4197;	// sequencer-master.scala:133:52, :185:52
      wire _T_4222 = io_op_bits_active_vfcmp ? _T_2304 & _T_9 | ~_T_9 & _T_4198 : _T_4198;	// sequencer-master.scala:133:52, :185:52
      wire _T_4223 = io_op_bits_active_vfcmp ? _T_2305 & _T_9 | ~_T_9 & _T_4199 : _T_4199;	// sequencer-master.scala:133:52, :185:52
      wire _T_4224 = io_op_bits_active_vfcmp ? _T_2306 & _T_9 | ~_T_9 & _T_4200 : _T_4200;	// sequencer-master.scala:133:52, :185:52
      wire _T_4225 = io_op_bits_active_vfconv ? _T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 & _T_4201 : _T_4201;	// sequencer-master.scala:131:52, :183:52
      wire _T_4226 = io_op_bits_active_vfconv ? _T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 & _T_4202 : _T_4202;	// sequencer-master.scala:131:52, :183:52
      wire _T_4227 = io_op_bits_active_vfconv ? _T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 & _T_4203 : _T_4203;	// sequencer-master.scala:131:52, :183:52
      wire _T_4228 = io_op_bits_active_vfconv ? _T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 & _T_4204 : _T_4204;	// sequencer-master.scala:131:52, :183:52
      wire _T_4229 = io_op_bits_active_vfconv ? _T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 & _T_4205 : _T_4205;	// sequencer-master.scala:131:52, :183:52
      wire _T_4230 = io_op_bits_active_vfconv ? _T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 & _T_4206 : _T_4206;	// sequencer-master.scala:131:52, :183:52
      wire _T_4231 = io_op_bits_active_vfconv ? _T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 & _T_4207 : _T_4207;	// sequencer-master.scala:131:52, :183:52
      wire _T_4232 = io_op_bits_active_vfconv ? _T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 & _T_4208 : _T_4208;	// sequencer-master.scala:131:52, :183:52
      wire _T_4233 = io_op_bits_active_vrpred ? _T_2238 & _T_9 | ~_T_9 & _T_4225 : _T_4225;	// sequencer-master.scala:131:52, :183:52
      wire _T_4234 = io_op_bits_active_vrpred ? _T_2242 & _T_9 | ~_T_9 & _T_4226 : _T_4226;	// sequencer-master.scala:131:52, :183:52
      wire _T_4235 = io_op_bits_active_vrpred ? _T_2246 & _T_9 | ~_T_9 & _T_4227 : _T_4227;	// sequencer-master.scala:131:52, :183:52
      wire _T_4236 = io_op_bits_active_vrpred ? _T_2250 & _T_9 | ~_T_9 & _T_4228 : _T_4228;	// sequencer-master.scala:131:52, :183:52
      wire _T_4237 = io_op_bits_active_vrpred ? _T_2254 & _T_9 | ~_T_9 & _T_4229 : _T_4229;	// sequencer-master.scala:131:52, :183:52
      wire _T_4238 = io_op_bits_active_vrpred ? _T_2258 & _T_9 | ~_T_9 & _T_4230 : _T_4230;	// sequencer-master.scala:131:52, :183:52
      wire _T_4239 = io_op_bits_active_vrpred ? _T_2262 & _T_9 | ~_T_9 & _T_4231 : _T_4231;	// sequencer-master.scala:131:52, :183:52
      wire _T_4240 = io_op_bits_active_vrpred ? _T_2266 & _T_9 | ~_T_9 & _T_4232 : _T_4232;	// sequencer-master.scala:131:52, :183:52
      wire _T_4241 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_9 | ~_T_9 & _T_4209 : _T_4209);	// sequencer-master.scala:132:52, :184:52
      wire _T_4242 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_9 | ~_T_9 & _T_4217 : _T_4217);	// sequencer-master.scala:133:52, :185:52
      wire _T_4243 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_9 | ~_T_9 & _T_4210 : _T_4210);	// sequencer-master.scala:132:52, :184:52
      wire _T_4244 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_9 | ~_T_9 & _T_4218 : _T_4218);	// sequencer-master.scala:133:52, :185:52
      wire _T_4245 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_9 | ~_T_9 & _T_4211 : _T_4211);	// sequencer-master.scala:132:52, :184:52
      wire _T_4246 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_9 | ~_T_9 & _T_4219 : _T_4219);	// sequencer-master.scala:133:52, :185:52
      wire _T_4247 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_9 | ~_T_9 & _T_4212 : _T_4212);	// sequencer-master.scala:132:52, :184:52
      wire _T_4248 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_9 | ~_T_9 & _T_4220 : _T_4220);	// sequencer-master.scala:133:52, :185:52
      wire _T_4249 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_9 | ~_T_9 & _T_4213 : _T_4213);	// sequencer-master.scala:132:52, :184:52
      wire _T_4250 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_9 | ~_T_9 & _T_4221 : _T_4221);	// sequencer-master.scala:133:52, :185:52
      wire _T_4251 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_9 | ~_T_9 & _T_4214 : _T_4214);	// sequencer-master.scala:132:52, :184:52
      wire _T_4252 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_9 | ~_T_9 & _T_4222 : _T_4222);	// sequencer-master.scala:133:52, :185:52
      wire _T_4253 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_9 | ~_T_9 & _T_4215 : _T_4215);	// sequencer-master.scala:132:52, :184:52
      wire _T_4254 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_9 | ~_T_9 & _T_4223 : _T_4223);	// sequencer-master.scala:133:52, :185:52
      wire _T_4255 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_9 | ~_T_9 & _T_4216 : _T_4216);	// sequencer-master.scala:132:52, :184:52
      wire _T_4256 = (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_9 | ~_T_9 & _T_4224 : _T_4224);	// sequencer-master.scala:133:52, :185:52
      wire _T_4257 = io_op_bits_active_vrfirst ? _T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 & _T_4233 : _T_4233;	// sequencer-master.scala:131:52, :183:52
      wire _T_4258 = io_op_bits_active_vrfirst ? _T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 & _T_4234 : _T_4234;	// sequencer-master.scala:131:52, :183:52
      wire _T_4259 = io_op_bits_active_vrfirst ? _T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 & _T_4235 : _T_4235;	// sequencer-master.scala:131:52, :183:52
      wire _T_4260 = io_op_bits_active_vrfirst ? _T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 & _T_4236 : _T_4236;	// sequencer-master.scala:131:52, :183:52
      wire _T_4261 = io_op_bits_active_vrfirst ? _T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 & _T_4237 : _T_4237;	// sequencer-master.scala:131:52, :183:52
      wire _T_4262 = io_op_bits_active_vrfirst ? _T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 & _T_4238 : _T_4238;	// sequencer-master.scala:131:52, :183:52
      wire _T_4263 = io_op_bits_active_vrfirst ? _T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 & _T_4239 : _T_4239;	// sequencer-master.scala:131:52, :183:52
      wire _T_4264 = io_op_bits_active_vrfirst ? _T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 & _T_4240 : _T_4240;	// sequencer-master.scala:131:52, :183:52
      wire _T_4265 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_132 | _T_2279 & _T_296 | _T_2238 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2269 & _T_9 | _T_2238 & _T_9 | ~_T_9 & _T_4257)) : _T_4257;	// sequencer-master.scala:131:52, :183:52
      wire _T_4266 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_133 | _T_2280 & _T_296 | _T_2242 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2270 & _T_9 | _T_2242 & _T_9 | ~_T_9 & _T_4258)) : _T_4258;	// sequencer-master.scala:131:52, :183:52
      wire _T_4267 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_134 | _T_2281 & _T_296 | _T_2246 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2271 & _T_9 | _T_2246 & _T_9 | ~_T_9 & _T_4259)) : _T_4259;	// sequencer-master.scala:131:52, :183:52
      wire _T_4268 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_135 | _T_2282 & _T_296 | _T_2250 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2272 & _T_9 | _T_2250 & _T_9 | ~_T_9 & _T_4260)) : _T_4260;	// sequencer-master.scala:131:52, :183:52
      wire _T_4269 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_136 | _T_2283 & _T_296 | _T_2254 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2273 & _T_9 | _T_2254 & _T_9 | ~_T_9 & _T_4261)) : _T_4261;	// sequencer-master.scala:131:52, :183:52
      wire _T_4270 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_137 | _T_2284 & _T_296 | _T_2258 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2274 & _T_9 | _T_2258 & _T_9 | ~_T_9 & _T_4262)) : _T_4262;	// sequencer-master.scala:131:52, :183:52
      wire _T_4271 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & _T_138 | _T_2285 & _T_296 | _T_2262 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2275 & _T_9 | _T_2262 & _T_9 | ~_T_9 & _T_4263)) : _T_4263;	// sequencer-master.scala:131:52, :183:52
      wire _T_4272 = io_op_bits_active_vamo ? ~_T_319 & (_T_296 & &_T_0 | _T_2286 & _T_296 | _T_2266 & _T_296 |
                ~_T_296 & ~_T_137 & (_T_2276 & _T_9 | _T_2266 & _T_9 | ~_T_9 & _T_4264)) : _T_4264;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4273 = io_op_bits_active_vamo ? _T_2308 & _T_319 | ~_T_319 & ~_T_296 & (_T_2308 & _T_137 | ~_T_137
                & ~_T_9 & _T_4241) : _T_4241;	// sequencer-master.scala:132:52, :184:52
      wire _T_4274 = io_op_bits_active_vamo ? _T_2309 & _T_319 | ~_T_319 & ~_T_296 & (_T_2309 & _T_137 | ~_T_137
                & ~_T_9 & _T_4243) : _T_4243;	// sequencer-master.scala:132:52, :184:52
      wire _T_4275 = io_op_bits_active_vamo ? _T_2310 & _T_319 | ~_T_319 & ~_T_296 & (_T_2310 & _T_137 | ~_T_137
                & ~_T_9 & _T_4245) : _T_4245;	// sequencer-master.scala:132:52, :184:52
      wire _T_4276 = io_op_bits_active_vamo ? _T_2311 & _T_319 | ~_T_319 & ~_T_296 & (_T_2311 & _T_137 | ~_T_137
                & ~_T_9 & _T_4247) : _T_4247;	// sequencer-master.scala:132:52, :184:52
      wire _T_4277 = io_op_bits_active_vamo ? _T_2312 & _T_319 | ~_T_319 & ~_T_296 & (_T_2312 & _T_137 | ~_T_137
                & ~_T_9 & _T_4249) : _T_4249;	// sequencer-master.scala:132:52, :184:52
      wire _T_4278 = io_op_bits_active_vamo ? _T_2313 & _T_319 | ~_T_319 & ~_T_296 & (_T_2313 & _T_137 | ~_T_137
                & ~_T_9 & _T_4251) : _T_4251;	// sequencer-master.scala:132:52, :184:52
      wire _T_4279 = io_op_bits_active_vamo ? _T_2314 & _T_319 | ~_T_319 & ~_T_296 & (_T_2314 & _T_137 | ~_T_137
                & ~_T_9 & _T_4253) : _T_4253;	// sequencer-master.scala:132:52, :184:52
      wire _T_4280 = io_op_bits_active_vamo ? _T_2315 & _T_319 | ~_T_319 & ~_T_296 & (_T_2315 & _T_137 | ~_T_137
                & ~_T_9 & _T_4255) : _T_4255;	// sequencer-master.scala:132:52, :184:52
      wire _T_4281 = io_op_bits_active_vamo ? _T_2299 & _T_319 | ~_T_319 & ~_T_296 & (_T_2299 & _T_137 | ~_T_137
                & ~_T_9 & _T_4242) : _T_4242;	// sequencer-master.scala:133:52, :185:52
      wire _T_4282 = io_op_bits_active_vamo ? _T_2300 & _T_319 | ~_T_319 & ~_T_296 & (_T_2300 & _T_137 | ~_T_137
                & ~_T_9 & _T_4244) : _T_4244;	// sequencer-master.scala:133:52, :185:52
      wire _T_4283 = io_op_bits_active_vamo ? _T_2301 & _T_319 | ~_T_319 & ~_T_296 & (_T_2301 & _T_137 | ~_T_137
                & ~_T_9 & _T_4246) : _T_4246;	// sequencer-master.scala:133:52, :185:52
      wire _T_4284 = io_op_bits_active_vamo ? _T_2302 & _T_319 | ~_T_319 & ~_T_296 & (_T_2302 & _T_137 | ~_T_137
                & ~_T_9 & _T_4248) : _T_4248;	// sequencer-master.scala:133:52, :185:52
      wire _T_4285 = io_op_bits_active_vamo ? _T_2303 & _T_319 | ~_T_319 & ~_T_296 & (_T_2303 & _T_137 | ~_T_137
                & ~_T_9 & _T_4250) : _T_4250;	// sequencer-master.scala:133:52, :185:52
      wire _T_4286 = io_op_bits_active_vamo ? _T_2304 & _T_319 | ~_T_319 & ~_T_296 & (_T_2304 & _T_137 | ~_T_137
                & ~_T_9 & _T_4252) : _T_4252;	// sequencer-master.scala:133:52, :185:52
      wire _T_4287 = io_op_bits_active_vamo ? _T_2305 & _T_319 | ~_T_319 & ~_T_296 & (_T_2305 & _T_137 | ~_T_137
                & ~_T_9 & _T_4254) : _T_4254;	// sequencer-master.scala:133:52, :185:52
      wire _T_4288 = io_op_bits_active_vamo ? _T_2306 & _T_319 | ~_T_319 & ~_T_296 & (_T_2306 & _T_137 | ~_T_137
                & ~_T_9 & _T_4256) : _T_4256;	// sequencer-master.scala:133:52, :185:52
      wire _T_4289 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2279 & _T_9 | _T_2238 & _T_9 | ~_T_9 &
                _T_4265) : _T_4265;	// sequencer-master.scala:131:52, :183:52
      wire _T_4290 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2280 & _T_9 | _T_2242 & _T_9 | ~_T_9 &
                _T_4266) : _T_4266;	// sequencer-master.scala:131:52, :183:52
      wire _T_4291 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2281 & _T_9 | _T_2246 & _T_9 | ~_T_9 &
                _T_4267) : _T_4267;	// sequencer-master.scala:131:52, :183:52
      wire _T_4292 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2282 & _T_9 | _T_2250 & _T_9 | ~_T_9 &
                _T_4268) : _T_4268;	// sequencer-master.scala:131:52, :183:52
      wire _T_4293 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2283 & _T_9 | _T_2254 & _T_9 | ~_T_9 &
                _T_4269) : _T_4269;	// sequencer-master.scala:131:52, :183:52
      wire _T_4294 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2284 & _T_9 | _T_2258 & _T_9 | ~_T_9 &
                _T_4270) : _T_4270;	// sequencer-master.scala:131:52, :183:52
      wire _T_4295 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2285 & _T_9 | _T_2262 & _T_9 | ~_T_9 &
                _T_4271) : _T_4271;	// sequencer-master.scala:131:52, :183:52
      wire _T_4296 = io_op_bits_active_vldx ? ~_T_296 & ~_T_137 & (_T_2286 & _T_9 | _T_2266 & _T_9 | ~_T_9 &
                _T_4272) : _T_4272;	// sequencer-master.scala:131:52, :183:52
      wire _T_4297 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2308 &
                _T_296 | ~_T_296 & (_T_2308 & _T_137 | ~_T_137 & ~_T_9 & _T_4273) : _T_4273);	// sequencer-master.scala:132:52, :184:52
      wire _T_4298 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2299 &
                _T_296 | ~_T_296 & (_T_2299 & _T_137 | ~_T_137 & ~_T_9 & _T_4281) : _T_4281);	// sequencer-master.scala:133:52, :185:52
      wire _T_4299 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2309 &
                _T_296 | ~_T_296 & (_T_2309 & _T_137 | ~_T_137 & ~_T_9 & _T_4274) : _T_4274);	// sequencer-master.scala:132:52, :184:52
      wire _T_4300 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2300 &
                _T_296 | ~_T_296 & (_T_2300 & _T_137 | ~_T_137 & ~_T_9 & _T_4282) : _T_4282);	// sequencer-master.scala:133:52, :185:52
      wire _T_4301 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2310 &
                _T_296 | ~_T_296 & (_T_2310 & _T_137 | ~_T_137 & ~_T_9 & _T_4275) : _T_4275);	// sequencer-master.scala:132:52, :184:52
      wire _T_4302 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2301 &
                _T_296 | ~_T_296 & (_T_2301 & _T_137 | ~_T_137 & ~_T_9 & _T_4283) : _T_4283);	// sequencer-master.scala:133:52, :185:52
      wire _T_4303 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2311 &
                _T_296 | ~_T_296 & (_T_2311 & _T_137 | ~_T_137 & ~_T_9 & _T_4276) : _T_4276);	// sequencer-master.scala:132:52, :184:52
      wire _T_4304 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2302 &
                _T_296 | ~_T_296 & (_T_2302 & _T_137 | ~_T_137 & ~_T_9 & _T_4284) : _T_4284);	// sequencer-master.scala:133:52, :185:52
      wire _T_4305 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2312 &
                _T_296 | ~_T_296 & (_T_2312 & _T_137 | ~_T_137 & ~_T_9 & _T_4277) : _T_4277);	// sequencer-master.scala:132:52, :184:52
      wire _T_4306 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2303 &
                _T_296 | ~_T_296 & (_T_2303 & _T_137 | ~_T_137 & ~_T_9 & _T_4285) : _T_4285);	// sequencer-master.scala:133:52, :185:52
      wire _T_4307 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2313 &
                _T_296 | ~_T_296 & (_T_2313 & _T_137 | ~_T_137 & ~_T_9 & _T_4278) : _T_4278);	// sequencer-master.scala:132:52, :184:52
      wire _T_4308 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2304 &
                _T_296 | ~_T_296 & (_T_2304 & _T_137 | ~_T_137 & ~_T_9 & _T_4286) : _T_4286);	// sequencer-master.scala:133:52, :185:52
      wire _T_4309 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2314 &
                _T_296 | ~_T_296 & (_T_2314 & _T_137 | ~_T_137 & ~_T_9 & _T_4279) : _T_4279);	// sequencer-master.scala:132:52, :184:52
      wire _T_4310 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2305 &
                _T_296 | ~_T_296 & (_T_2305 & _T_137 | ~_T_137 & ~_T_9 & _T_4287) : _T_4287);	// sequencer-master.scala:133:52, :185:52
      wire _T_4311 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2315 &
                _T_296 | ~_T_296 & (_T_2315 & _T_137 | ~_T_137 & ~_T_9 & _T_4280) : _T_4280);	// sequencer-master.scala:132:52, :184:52
      wire _T_4312 = (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vldx ? _T_2306 &
                _T_296 | ~_T_296 & (_T_2306 & _T_137 | ~_T_137 & ~_T_9 & _T_4288) : _T_4288);	// sequencer-master.scala:133:52, :185:52
      wire _T_4313 = io_op_bits_active_vstx ? _T_296 & _T_132 | _T_2299 & _T_296 | _T_2238 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2279 & _T_9 | _T_2238 & _T_9 | ~_T_9 & _T_4289) : _T_4289;	// sequencer-master.scala:131:52, :183:52
      wire _T_4314 = io_op_bits_active_vstx ? _T_296 & _T_133 | _T_2300 & _T_296 | _T_2242 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2280 & _T_9 | _T_2242 & _T_9 | ~_T_9 & _T_4290) : _T_4290;	// sequencer-master.scala:131:52, :183:52
      wire _T_4315 = io_op_bits_active_vstx ? _T_296 & _T_134 | _T_2301 & _T_296 | _T_2246 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2281 & _T_9 | _T_2246 & _T_9 | ~_T_9 & _T_4291) : _T_4291;	// sequencer-master.scala:131:52, :183:52
      wire _T_4316 = io_op_bits_active_vstx ? _T_296 & _T_135 | _T_2302 & _T_296 | _T_2250 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2282 & _T_9 | _T_2250 & _T_9 | ~_T_9 & _T_4292) : _T_4292;	// sequencer-master.scala:131:52, :183:52
      wire _T_4317 = io_op_bits_active_vstx ? _T_296 & _T_136 | _T_2303 & _T_296 | _T_2254 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2283 & _T_9 | _T_2254 & _T_9 | ~_T_9 & _T_4293) : _T_4293;	// sequencer-master.scala:131:52, :183:52
      wire _T_4318 = io_op_bits_active_vstx ? _T_296 & _T_137 | _T_2304 & _T_296 | _T_2258 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2284 & _T_9 | _T_2258 & _T_9 | ~_T_9 & _T_4294) : _T_4294;	// sequencer-master.scala:131:52, :183:52
      wire _T_4319 = io_op_bits_active_vstx ? _T_296 & _T_138 | _T_2305 & _T_296 | _T_2262 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2285 & _T_9 | _T_2262 & _T_9 | ~_T_9 & _T_4295) : _T_4295;	// sequencer-master.scala:131:52, :183:52
      wire _T_4320 = io_op_bits_active_vstx ? _T_296 & &_T_0 | _T_2306 & _T_296 | _T_2266 & _T_296 | ~_T_296 &
                ~_T_137 & (_T_2286 & _T_9 | _T_2266 & _T_9 | ~_T_9 & _T_4296) : _T_4296;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4321 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2238 & _T_9 | ~_T_9 & _T_4313) : _T_4313;	// sequencer-master.scala:131:52, :183:52
      wire _T_4322 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2242 & _T_9 | ~_T_9 & _T_4314) : _T_4314;	// sequencer-master.scala:131:52, :183:52
      wire _T_4323 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2246 & _T_9 | ~_T_9 & _T_4315) : _T_4315;	// sequencer-master.scala:131:52, :183:52
      wire _T_4324 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2250 & _T_9 | ~_T_9 & _T_4316) : _T_4316;	// sequencer-master.scala:131:52, :183:52
      wire _T_4325 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2254 & _T_9 | ~_T_9 & _T_4317) : _T_4317;	// sequencer-master.scala:131:52, :183:52
      wire _T_4326 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2258 & _T_9 | ~_T_9 & _T_4318) : _T_4318;	// sequencer-master.scala:131:52, :183:52
      wire _T_4327 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2262 & _T_9 | ~_T_9 & _T_4319) : _T_4319;	// sequencer-master.scala:131:52, :183:52
      wire _T_4328 = io_op_bits_active_vld ? ~_T_296 & ~_T_137 & (_T_2266 & _T_9 | ~_T_9 & _T_4320) : _T_4320;	// sequencer-master.scala:131:52, :183:52
      wire _T_4329 = io_op_bits_active_vint ? _T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 &
                e_6_raw_0 : e_6_raw_0;	// sequencer-master.scala:131:52, :183:52
      wire _T_4330 = io_op_bits_active_vint ? _T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 &
                e_6_raw_1 : e_6_raw_1;	// sequencer-master.scala:131:52, :183:52
      wire _T_4331 = io_op_bits_active_vint ? _T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 &
                e_6_raw_2 : e_6_raw_2;	// sequencer-master.scala:131:52, :183:52
      wire _T_4332 = io_op_bits_active_vint ? _T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 &
                e_6_raw_3 : e_6_raw_3;	// sequencer-master.scala:131:52, :183:52
      wire _T_4333 = io_op_bits_active_vint ? _T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 &
                e_6_raw_4 : e_6_raw_4;	// sequencer-master.scala:131:52, :183:52
      wire _T_4334 = io_op_bits_active_vint ? _T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 &
                e_6_raw_5 : e_6_raw_5;	// sequencer-master.scala:131:52, :183:52
      wire _T_4335 = io_op_bits_active_vint ? _T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 &
                e_6_raw_6 : e_6_raw_6;	// sequencer-master.scala:131:52, :183:52
      wire _T_4336 = io_op_bits_active_vint ? _T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 &
                e_6_raw_7 : e_6_raw_7;	// sequencer-master.scala:131:52, :183:52
      wire _T_4337 = io_op_bits_active_vint ? _T_2308 & _T_10 | ~_T_10 & e_6_war_0 : e_6_war_0;	// sequencer-master.scala:132:52, :184:52
      wire _T_4338 = io_op_bits_active_vint ? _T_2309 & _T_10 | ~_T_10 & e_6_war_1 : e_6_war_1;	// sequencer-master.scala:132:52, :184:52
      wire _T_4339 = io_op_bits_active_vint ? _T_2310 & _T_10 | ~_T_10 & e_6_war_2 : e_6_war_2;	// sequencer-master.scala:132:52, :184:52
      wire _T_4340 = io_op_bits_active_vint ? _T_2311 & _T_10 | ~_T_10 & e_6_war_3 : e_6_war_3;	// sequencer-master.scala:132:52, :184:52
      wire _T_4341 = io_op_bits_active_vint ? _T_2312 & _T_10 | ~_T_10 & e_6_war_4 : e_6_war_4;	// sequencer-master.scala:132:52, :184:52
      wire _T_4342 = io_op_bits_active_vint ? _T_2313 & _T_10 | ~_T_10 & e_6_war_5 : e_6_war_5;	// sequencer-master.scala:132:52, :184:52
      wire _T_4343 = io_op_bits_active_vint ? _T_2314 & _T_10 | ~_T_10 & e_6_war_6 : e_6_war_6;	// sequencer-master.scala:132:52, :184:52
      wire _T_4344 = io_op_bits_active_vint ? _T_2315 & _T_10 | ~_T_10 & e_6_war_7 : e_6_war_7;	// sequencer-master.scala:132:52, :184:52
      wire _T_4345 = io_op_bits_active_vint ? _T_2299 & _T_10 | ~_T_10 & e_6_waw_0 : e_6_waw_0;	// sequencer-master.scala:133:52, :185:52
      wire _T_4346 = io_op_bits_active_vint ? _T_2300 & _T_10 | ~_T_10 & e_6_waw_1 : e_6_waw_1;	// sequencer-master.scala:133:52, :185:52
      wire _T_4347 = io_op_bits_active_vint ? _T_2301 & _T_10 | ~_T_10 & e_6_waw_2 : e_6_waw_2;	// sequencer-master.scala:133:52, :185:52
      wire _T_4348 = io_op_bits_active_vint ? _T_2302 & _T_10 | ~_T_10 & e_6_waw_3 : e_6_waw_3;	// sequencer-master.scala:133:52, :185:52
      wire _T_4349 = io_op_bits_active_vint ? _T_2303 & _T_10 | ~_T_10 & e_6_waw_4 : e_6_waw_4;	// sequencer-master.scala:133:52, :185:52
      wire _T_4350 = io_op_bits_active_vint ? _T_2304 & _T_10 | ~_T_10 & e_6_waw_5 : e_6_waw_5;	// sequencer-master.scala:133:52, :185:52
      wire _T_4351 = io_op_bits_active_vint ? _T_2305 & _T_10 | ~_T_10 & e_6_waw_6 : e_6_waw_6;	// sequencer-master.scala:133:52, :185:52
      wire _T_4352 = io_op_bits_active_vint ? _T_2306 & _T_10 | ~_T_10 & e_6_waw_7 : e_6_waw_7;	// sequencer-master.scala:133:52, :185:52
      wire _T_4353 = io_op_bits_active_vipred ? _T_2289 & _T_10 | _T_2279 & _T_10 | _T_2269 & _T_10 | ~_T_10 &
                _T_4329 : _T_4329;	// sequencer-master.scala:131:52, :183:52
      wire _T_4354 = io_op_bits_active_vipred ? _T_2290 & _T_10 | _T_2280 & _T_10 | _T_2270 & _T_10 | ~_T_10 &
                _T_4330 : _T_4330;	// sequencer-master.scala:131:52, :183:52
      wire _T_4355 = io_op_bits_active_vipred ? _T_2291 & _T_10 | _T_2281 & _T_10 | _T_2271 & _T_10 | ~_T_10 &
                _T_4331 : _T_4331;	// sequencer-master.scala:131:52, :183:52
      wire _T_4356 = io_op_bits_active_vipred ? _T_2292 & _T_10 | _T_2282 & _T_10 | _T_2272 & _T_10 | ~_T_10 &
                _T_4332 : _T_4332;	// sequencer-master.scala:131:52, :183:52
      wire _T_4357 = io_op_bits_active_vipred ? _T_2293 & _T_10 | _T_2283 & _T_10 | _T_2273 & _T_10 | ~_T_10 &
                _T_4333 : _T_4333;	// sequencer-master.scala:131:52, :183:52
      wire _T_4358 = io_op_bits_active_vipred ? _T_2294 & _T_10 | _T_2284 & _T_10 | _T_2274 & _T_10 | ~_T_10 &
                _T_4334 : _T_4334;	// sequencer-master.scala:131:52, :183:52
      wire _T_4359 = io_op_bits_active_vipred ? _T_2295 & _T_10 | _T_2285 & _T_10 | _T_2275 & _T_10 | ~_T_10 &
                _T_4335 : _T_4335;	// sequencer-master.scala:131:52, :183:52
      wire _T_4360 = io_op_bits_active_vipred ? _T_2296 & _T_10 | _T_2286 & _T_10 | _T_2276 & _T_10 | ~_T_10 &
                _T_4336 : _T_4336;	// sequencer-master.scala:131:52, :183:52
      wire _T_4361 = io_op_bits_active_vipred ? _T_2308 & _T_10 | ~_T_10 & _T_4337 : _T_4337;	// sequencer-master.scala:132:52, :184:52
      wire _T_4362 = io_op_bits_active_vipred ? _T_2309 & _T_10 | ~_T_10 & _T_4338 : _T_4338;	// sequencer-master.scala:132:52, :184:52
      wire _T_4363 = io_op_bits_active_vipred ? _T_2310 & _T_10 | ~_T_10 & _T_4339 : _T_4339;	// sequencer-master.scala:132:52, :184:52
      wire _T_4364 = io_op_bits_active_vipred ? _T_2311 & _T_10 | ~_T_10 & _T_4340 : _T_4340;	// sequencer-master.scala:132:52, :184:52
      wire _T_4365 = io_op_bits_active_vipred ? _T_2312 & _T_10 | ~_T_10 & _T_4341 : _T_4341;	// sequencer-master.scala:132:52, :184:52
      wire _T_4366 = io_op_bits_active_vipred ? _T_2313 & _T_10 | ~_T_10 & _T_4342 : _T_4342;	// sequencer-master.scala:132:52, :184:52
      wire _T_4367 = io_op_bits_active_vipred ? _T_2314 & _T_10 | ~_T_10 & _T_4343 : _T_4343;	// sequencer-master.scala:132:52, :184:52
      wire _T_4368 = io_op_bits_active_vipred ? _T_2315 & _T_10 | ~_T_10 & _T_4344 : _T_4344;	// sequencer-master.scala:132:52, :184:52
      wire _T_4369 = io_op_bits_active_vipred ? _T_2299 & _T_10 | ~_T_10 & _T_4345 : _T_4345;	// sequencer-master.scala:133:52, :185:52
      wire _T_4370 = io_op_bits_active_vipred ? _T_2300 & _T_10 | ~_T_10 & _T_4346 : _T_4346;	// sequencer-master.scala:133:52, :185:52
      wire _T_4371 = io_op_bits_active_vipred ? _T_2301 & _T_10 | ~_T_10 & _T_4347 : _T_4347;	// sequencer-master.scala:133:52, :185:52
      wire _T_4372 = io_op_bits_active_vipred ? _T_2302 & _T_10 | ~_T_10 & _T_4348 : _T_4348;	// sequencer-master.scala:133:52, :185:52
      wire _T_4373 = io_op_bits_active_vipred ? _T_2303 & _T_10 | ~_T_10 & _T_4349 : _T_4349;	// sequencer-master.scala:133:52, :185:52
      wire _T_4374 = io_op_bits_active_vipred ? _T_2304 & _T_10 | ~_T_10 & _T_4350 : _T_4350;	// sequencer-master.scala:133:52, :185:52
      wire _T_4375 = io_op_bits_active_vipred ? _T_2305 & _T_10 | ~_T_10 & _T_4351 : _T_4351;	// sequencer-master.scala:133:52, :185:52
      wire _T_4376 = io_op_bits_active_vipred ? _T_2306 & _T_10 | ~_T_10 & _T_4352 : _T_4352;	// sequencer-master.scala:133:52, :185:52
      wire _T_4377 = io_op_bits_active_vimul ? _T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 &
                _T_4353 : _T_4353;	// sequencer-master.scala:131:52, :183:52
      wire _T_4378 = io_op_bits_active_vimul ? _T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 &
                _T_4354 : _T_4354;	// sequencer-master.scala:131:52, :183:52
      wire _T_4379 = io_op_bits_active_vimul ? _T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 &
                _T_4355 : _T_4355;	// sequencer-master.scala:131:52, :183:52
      wire _T_4380 = io_op_bits_active_vimul ? _T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 &
                _T_4356 : _T_4356;	// sequencer-master.scala:131:52, :183:52
      wire _T_4381 = io_op_bits_active_vimul ? _T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 &
                _T_4357 : _T_4357;	// sequencer-master.scala:131:52, :183:52
      wire _T_4382 = io_op_bits_active_vimul ? _T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 &
                _T_4358 : _T_4358;	// sequencer-master.scala:131:52, :183:52
      wire _T_4383 = io_op_bits_active_vimul ? _T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 &
                _T_4359 : _T_4359;	// sequencer-master.scala:131:52, :183:52
      wire _T_4384 = io_op_bits_active_vimul ? _T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 &
                _T_4360 : _T_4360;	// sequencer-master.scala:131:52, :183:52
      wire _T_4385 = io_op_bits_active_vimul ? _T_2308 & _T_10 | ~_T_10 & _T_4361 : _T_4361;	// sequencer-master.scala:132:52, :184:52
      wire _T_4386 = io_op_bits_active_vimul ? _T_2309 & _T_10 | ~_T_10 & _T_4362 : _T_4362;	// sequencer-master.scala:132:52, :184:52
      wire _T_4387 = io_op_bits_active_vimul ? _T_2310 & _T_10 | ~_T_10 & _T_4363 : _T_4363;	// sequencer-master.scala:132:52, :184:52
      wire _T_4388 = io_op_bits_active_vimul ? _T_2311 & _T_10 | ~_T_10 & _T_4364 : _T_4364;	// sequencer-master.scala:132:52, :184:52
      wire _T_4389 = io_op_bits_active_vimul ? _T_2312 & _T_10 | ~_T_10 & _T_4365 : _T_4365;	// sequencer-master.scala:132:52, :184:52
      wire _T_4390 = io_op_bits_active_vimul ? _T_2313 & _T_10 | ~_T_10 & _T_4366 : _T_4366;	// sequencer-master.scala:132:52, :184:52
      wire _T_4391 = io_op_bits_active_vimul ? _T_2314 & _T_10 | ~_T_10 & _T_4367 : _T_4367;	// sequencer-master.scala:132:52, :184:52
      wire _T_4392 = io_op_bits_active_vimul ? _T_2315 & _T_10 | ~_T_10 & _T_4368 : _T_4368;	// sequencer-master.scala:132:52, :184:52
      wire _T_4393 = io_op_bits_active_vimul ? _T_2299 & _T_10 | ~_T_10 & _T_4369 : _T_4369;	// sequencer-master.scala:133:52, :185:52
      wire _T_4394 = io_op_bits_active_vimul ? _T_2300 & _T_10 | ~_T_10 & _T_4370 : _T_4370;	// sequencer-master.scala:133:52, :185:52
      wire _T_4395 = io_op_bits_active_vimul ? _T_2301 & _T_10 | ~_T_10 & _T_4371 : _T_4371;	// sequencer-master.scala:133:52, :185:52
      wire _T_4396 = io_op_bits_active_vimul ? _T_2302 & _T_10 | ~_T_10 & _T_4372 : _T_4372;	// sequencer-master.scala:133:52, :185:52
      wire _T_4397 = io_op_bits_active_vimul ? _T_2303 & _T_10 | ~_T_10 & _T_4373 : _T_4373;	// sequencer-master.scala:133:52, :185:52
      wire _T_4398 = io_op_bits_active_vimul ? _T_2304 & _T_10 | ~_T_10 & _T_4374 : _T_4374;	// sequencer-master.scala:133:52, :185:52
      wire _T_4399 = io_op_bits_active_vimul ? _T_2305 & _T_10 | ~_T_10 & _T_4375 : _T_4375;	// sequencer-master.scala:133:52, :185:52
      wire _T_4400 = io_op_bits_active_vimul ? _T_2306 & _T_10 | ~_T_10 & _T_4376 : _T_4376;	// sequencer-master.scala:133:52, :185:52
      wire _T_4401 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 & _T_10 |
                ~_T_10 & _T_4377) : _T_4377;	// sequencer-master.scala:131:52, :183:52
      wire _T_4402 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 & _T_10 |
                ~_T_10 & _T_4378) : _T_4378;	// sequencer-master.scala:131:52, :183:52
      wire _T_4403 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 & _T_10 |
                ~_T_10 & _T_4379) : _T_4379;	// sequencer-master.scala:131:52, :183:52
      wire _T_4404 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 & _T_10 |
                ~_T_10 & _T_4380) : _T_4380;	// sequencer-master.scala:131:52, :183:52
      wire _T_4405 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 & _T_10 |
                ~_T_10 & _T_4381) : _T_4381;	// sequencer-master.scala:131:52, :183:52
      wire _T_4406 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 & _T_10 |
                ~_T_10 & _T_4382) : _T_4382;	// sequencer-master.scala:131:52, :183:52
      wire _T_4407 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 & _T_10 |
                ~_T_10 & _T_4383) : _T_4383;	// sequencer-master.scala:131:52, :183:52
      wire _T_4408 = io_op_bits_active_vidiv ? ~_T_138 & (_T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 & _T_10 |
                ~_T_10 & _T_4384) : _T_4384;	// sequencer-master.scala:131:52, :183:52
      wire _T_4409 = io_op_bits_active_vidiv ? _T_2308 & _T_138 | ~_T_138 & (_T_2308 & _T_10 | ~_T_10 & _T_4385)
                : _T_4385;	// sequencer-master.scala:132:52, :184:52
      wire _T_4410 = io_op_bits_active_vidiv ? _T_2309 & _T_138 | ~_T_138 & (_T_2309 & _T_10 | ~_T_10 & _T_4386)
                : _T_4386;	// sequencer-master.scala:132:52, :184:52
      wire _T_4411 = io_op_bits_active_vidiv ? _T_2310 & _T_138 | ~_T_138 & (_T_2310 & _T_10 | ~_T_10 & _T_4387)
                : _T_4387;	// sequencer-master.scala:132:52, :184:52
      wire _T_4412 = io_op_bits_active_vidiv ? _T_2311 & _T_138 | ~_T_138 & (_T_2311 & _T_10 | ~_T_10 & _T_4388)
                : _T_4388;	// sequencer-master.scala:132:52, :184:52
      wire _T_4413 = io_op_bits_active_vidiv ? _T_2312 & _T_138 | ~_T_138 & (_T_2312 & _T_10 | ~_T_10 & _T_4389)
                : _T_4389;	// sequencer-master.scala:132:52, :184:52
      wire _T_4414 = io_op_bits_active_vidiv ? _T_2313 & _T_138 | ~_T_138 & (_T_2313 & _T_10 | ~_T_10 & _T_4390)
                : _T_4390;	// sequencer-master.scala:132:52, :184:52
      wire _T_4415 = io_op_bits_active_vidiv ? _T_2314 & _T_138 | ~_T_138 & (_T_2314 & _T_10 | ~_T_10 & _T_4391)
                : _T_4391;	// sequencer-master.scala:132:52, :184:52
      wire _T_4416 = io_op_bits_active_vidiv ? _T_2315 & _T_138 | ~_T_138 & (_T_2315 & _T_10 | ~_T_10 & _T_4392)
                : _T_4392;	// sequencer-master.scala:132:52, :184:52
      wire _T_4417 = io_op_bits_active_vidiv ? _T_2299 & _T_138 | ~_T_138 & (_T_2299 & _T_10 | ~_T_10 & _T_4393)
                : _T_4393;	// sequencer-master.scala:133:52, :185:52
      wire _T_4418 = io_op_bits_active_vidiv ? _T_2300 & _T_138 | ~_T_138 & (_T_2300 & _T_10 | ~_T_10 & _T_4394)
                : _T_4394;	// sequencer-master.scala:133:52, :185:52
      wire _T_4419 = io_op_bits_active_vidiv ? _T_2301 & _T_138 | ~_T_138 & (_T_2301 & _T_10 | ~_T_10 & _T_4395)
                : _T_4395;	// sequencer-master.scala:133:52, :185:52
      wire _T_4420 = io_op_bits_active_vidiv ? _T_2302 & _T_138 | ~_T_138 & (_T_2302 & _T_10 | ~_T_10 & _T_4396)
                : _T_4396;	// sequencer-master.scala:133:52, :185:52
      wire _T_4421 = io_op_bits_active_vidiv ? _T_2303 & _T_138 | ~_T_138 & (_T_2303 & _T_10 | ~_T_10 & _T_4397)
                : _T_4397;	// sequencer-master.scala:133:52, :185:52
      wire _T_4422 = io_op_bits_active_vidiv ? _T_2304 & _T_138 | ~_T_138 & (_T_2304 & _T_10 | ~_T_10 & _T_4398)
                : _T_4398;	// sequencer-master.scala:133:52, :185:52
      wire _T_4423 = io_op_bits_active_vidiv ? _T_2305 & _T_138 | ~_T_138 & (_T_2305 & _T_10 | ~_T_10 & _T_4399)
                : _T_4399;	// sequencer-master.scala:133:52, :185:52
      wire _T_4424 = io_op_bits_active_vidiv ? _T_2306 & _T_138 | ~_T_138 & (_T_2306 & _T_10 | ~_T_10 & _T_4400)
                : _T_4400;	// sequencer-master.scala:133:52, :185:52
      wire _T_4425 = io_op_bits_active_vfma ? _T_2289 & _T_10 | _T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 &
                _T_10 | ~_T_10 & _T_4401 : _T_4401;	// sequencer-master.scala:131:52, :183:52
      wire _T_4426 = io_op_bits_active_vfma ? _T_2290 & _T_10 | _T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 &
                _T_10 | ~_T_10 & _T_4402 : _T_4402;	// sequencer-master.scala:131:52, :183:52
      wire _T_4427 = io_op_bits_active_vfma ? _T_2291 & _T_10 | _T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 &
                _T_10 | ~_T_10 & _T_4403 : _T_4403;	// sequencer-master.scala:131:52, :183:52
      wire _T_4428 = io_op_bits_active_vfma ? _T_2292 & _T_10 | _T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 &
                _T_10 | ~_T_10 & _T_4404 : _T_4404;	// sequencer-master.scala:131:52, :183:52
      wire _T_4429 = io_op_bits_active_vfma ? _T_2293 & _T_10 | _T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 &
                _T_10 | ~_T_10 & _T_4405 : _T_4405;	// sequencer-master.scala:131:52, :183:52
      wire _T_4430 = io_op_bits_active_vfma ? _T_2294 & _T_10 | _T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 &
                _T_10 | ~_T_10 & _T_4406 : _T_4406;	// sequencer-master.scala:131:52, :183:52
      wire _T_4431 = io_op_bits_active_vfma ? _T_2295 & _T_10 | _T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 &
                _T_10 | ~_T_10 & _T_4407 : _T_4407;	// sequencer-master.scala:131:52, :183:52
      wire _T_4432 = io_op_bits_active_vfma ? _T_2296 & _T_10 | _T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 &
                _T_10 | ~_T_10 & _T_4408 : _T_4408;	// sequencer-master.scala:131:52, :183:52
      wire _T_4433 = io_op_bits_active_vfma ? _T_2308 & _T_10 | ~_T_10 & _T_4409 : _T_4409;	// sequencer-master.scala:132:52, :184:52
      wire _T_4434 = io_op_bits_active_vfma ? _T_2309 & _T_10 | ~_T_10 & _T_4410 : _T_4410;	// sequencer-master.scala:132:52, :184:52
      wire _T_4435 = io_op_bits_active_vfma ? _T_2310 & _T_10 | ~_T_10 & _T_4411 : _T_4411;	// sequencer-master.scala:132:52, :184:52
      wire _T_4436 = io_op_bits_active_vfma ? _T_2311 & _T_10 | ~_T_10 & _T_4412 : _T_4412;	// sequencer-master.scala:132:52, :184:52
      wire _T_4437 = io_op_bits_active_vfma ? _T_2312 & _T_10 | ~_T_10 & _T_4413 : _T_4413;	// sequencer-master.scala:132:52, :184:52
      wire _T_4438 = io_op_bits_active_vfma ? _T_2313 & _T_10 | ~_T_10 & _T_4414 : _T_4414;	// sequencer-master.scala:132:52, :184:52
      wire _T_4439 = io_op_bits_active_vfma ? _T_2314 & _T_10 | ~_T_10 & _T_4415 : _T_4415;	// sequencer-master.scala:132:52, :184:52
      wire _T_4440 = io_op_bits_active_vfma ? _T_2315 & _T_10 | ~_T_10 & _T_4416 : _T_4416;	// sequencer-master.scala:132:52, :184:52
      wire _T_4441 = io_op_bits_active_vfma ? _T_2299 & _T_10 | ~_T_10 & _T_4417 : _T_4417;	// sequencer-master.scala:133:52, :185:52
      wire _T_4442 = io_op_bits_active_vfma ? _T_2300 & _T_10 | ~_T_10 & _T_4418 : _T_4418;	// sequencer-master.scala:133:52, :185:52
      wire _T_4443 = io_op_bits_active_vfma ? _T_2301 & _T_10 | ~_T_10 & _T_4419 : _T_4419;	// sequencer-master.scala:133:52, :185:52
      wire _T_4444 = io_op_bits_active_vfma ? _T_2302 & _T_10 | ~_T_10 & _T_4420 : _T_4420;	// sequencer-master.scala:133:52, :185:52
      wire _T_4445 = io_op_bits_active_vfma ? _T_2303 & _T_10 | ~_T_10 & _T_4421 : _T_4421;	// sequencer-master.scala:133:52, :185:52
      wire _T_4446 = io_op_bits_active_vfma ? _T_2304 & _T_10 | ~_T_10 & _T_4422 : _T_4422;	// sequencer-master.scala:133:52, :185:52
      wire _T_4447 = io_op_bits_active_vfma ? _T_2305 & _T_10 | ~_T_10 & _T_4423 : _T_4423;	// sequencer-master.scala:133:52, :185:52
      wire _T_4448 = io_op_bits_active_vfma ? _T_2306 & _T_10 | ~_T_10 & _T_4424 : _T_4424;	// sequencer-master.scala:133:52, :185:52
      wire _T_4449 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 & _T_10 |
                ~_T_10 & _T_4425) : _T_4425;	// sequencer-master.scala:131:52, :183:52
      wire _T_4450 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 & _T_10 |
                ~_T_10 & _T_4426) : _T_4426;	// sequencer-master.scala:131:52, :183:52
      wire _T_4451 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 & _T_10 |
                ~_T_10 & _T_4427) : _T_4427;	// sequencer-master.scala:131:52, :183:52
      wire _T_4452 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 & _T_10 |
                ~_T_10 & _T_4428) : _T_4428;	// sequencer-master.scala:131:52, :183:52
      wire _T_4453 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 & _T_10 |
                ~_T_10 & _T_4429) : _T_4429;	// sequencer-master.scala:131:52, :183:52
      wire _T_4454 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 & _T_10 |
                ~_T_10 & _T_4430) : _T_4430;	// sequencer-master.scala:131:52, :183:52
      wire _T_4455 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 & _T_10 |
                ~_T_10 & _T_4431) : _T_4431;	// sequencer-master.scala:131:52, :183:52
      wire _T_4456 = io_op_bits_active_vfdiv ? ~_T_138 & (_T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 & _T_10 |
                ~_T_10 & _T_4432) : _T_4432;	// sequencer-master.scala:131:52, :183:52
      wire _T_4457 = io_op_bits_active_vfdiv ? _T_2308 & _T_138 | ~_T_138 & (_T_2308 & _T_10 | ~_T_10 & _T_4433)
                : _T_4433;	// sequencer-master.scala:132:52, :184:52
      wire _T_4458 = io_op_bits_active_vfdiv ? _T_2309 & _T_138 | ~_T_138 & (_T_2309 & _T_10 | ~_T_10 & _T_4434)
                : _T_4434;	// sequencer-master.scala:132:52, :184:52
      wire _T_4459 = io_op_bits_active_vfdiv ? _T_2310 & _T_138 | ~_T_138 & (_T_2310 & _T_10 | ~_T_10 & _T_4435)
                : _T_4435;	// sequencer-master.scala:132:52, :184:52
      wire _T_4460 = io_op_bits_active_vfdiv ? _T_2311 & _T_138 | ~_T_138 & (_T_2311 & _T_10 | ~_T_10 & _T_4436)
                : _T_4436;	// sequencer-master.scala:132:52, :184:52
      wire _T_4461 = io_op_bits_active_vfdiv ? _T_2312 & _T_138 | ~_T_138 & (_T_2312 & _T_10 | ~_T_10 & _T_4437)
                : _T_4437;	// sequencer-master.scala:132:52, :184:52
      wire _T_4462 = io_op_bits_active_vfdiv ? _T_2313 & _T_138 | ~_T_138 & (_T_2313 & _T_10 | ~_T_10 & _T_4438)
                : _T_4438;	// sequencer-master.scala:132:52, :184:52
      wire _T_4463 = io_op_bits_active_vfdiv ? _T_2314 & _T_138 | ~_T_138 & (_T_2314 & _T_10 | ~_T_10 & _T_4439)
                : _T_4439;	// sequencer-master.scala:132:52, :184:52
      wire _T_4464 = io_op_bits_active_vfdiv ? _T_2315 & _T_138 | ~_T_138 & (_T_2315 & _T_10 | ~_T_10 & _T_4440)
                : _T_4440;	// sequencer-master.scala:132:52, :184:52
      wire _T_4465 = io_op_bits_active_vfdiv ? _T_2299 & _T_138 | ~_T_138 & (_T_2299 & _T_10 | ~_T_10 & _T_4441)
                : _T_4441;	// sequencer-master.scala:133:52, :185:52
      wire _T_4466 = io_op_bits_active_vfdiv ? _T_2300 & _T_138 | ~_T_138 & (_T_2300 & _T_10 | ~_T_10 & _T_4442)
                : _T_4442;	// sequencer-master.scala:133:52, :185:52
      wire _T_4467 = io_op_bits_active_vfdiv ? _T_2301 & _T_138 | ~_T_138 & (_T_2301 & _T_10 | ~_T_10 & _T_4443)
                : _T_4443;	// sequencer-master.scala:133:52, :185:52
      wire _T_4468 = io_op_bits_active_vfdiv ? _T_2302 & _T_138 | ~_T_138 & (_T_2302 & _T_10 | ~_T_10 & _T_4444)
                : _T_4444;	// sequencer-master.scala:133:52, :185:52
      wire _T_4469 = io_op_bits_active_vfdiv ? _T_2303 & _T_138 | ~_T_138 & (_T_2303 & _T_10 | ~_T_10 & _T_4445)
                : _T_4445;	// sequencer-master.scala:133:52, :185:52
      wire _T_4470 = io_op_bits_active_vfdiv ? _T_2304 & _T_138 | ~_T_138 & (_T_2304 & _T_10 | ~_T_10 & _T_4446)
                : _T_4446;	// sequencer-master.scala:133:52, :185:52
      wire _T_4471 = io_op_bits_active_vfdiv ? _T_2305 & _T_138 | ~_T_138 & (_T_2305 & _T_10 | ~_T_10 & _T_4447)
                : _T_4447;	// sequencer-master.scala:133:52, :185:52
      wire _T_4472 = io_op_bits_active_vfdiv ? _T_2306 & _T_138 | ~_T_138 & (_T_2306 & _T_10 | ~_T_10 & _T_4448)
                : _T_4448;	// sequencer-master.scala:133:52, :185:52
      wire _T_4473 = io_op_bits_active_vfcmp ? _T_2279 & _T_10 | _T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 &
                _T_4449 : _T_4449;	// sequencer-master.scala:131:52, :183:52
      wire _T_4474 = io_op_bits_active_vfcmp ? _T_2280 & _T_10 | _T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 &
                _T_4450 : _T_4450;	// sequencer-master.scala:131:52, :183:52
      wire _T_4475 = io_op_bits_active_vfcmp ? _T_2281 & _T_10 | _T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 &
                _T_4451 : _T_4451;	// sequencer-master.scala:131:52, :183:52
      wire _T_4476 = io_op_bits_active_vfcmp ? _T_2282 & _T_10 | _T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 &
                _T_4452 : _T_4452;	// sequencer-master.scala:131:52, :183:52
      wire _T_4477 = io_op_bits_active_vfcmp ? _T_2283 & _T_10 | _T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 &
                _T_4453 : _T_4453;	// sequencer-master.scala:131:52, :183:52
      wire _T_4478 = io_op_bits_active_vfcmp ? _T_2284 & _T_10 | _T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 &
                _T_4454 : _T_4454;	// sequencer-master.scala:131:52, :183:52
      wire _T_4479 = io_op_bits_active_vfcmp ? _T_2285 & _T_10 | _T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 &
                _T_4455 : _T_4455;	// sequencer-master.scala:131:52, :183:52
      wire _T_4480 = io_op_bits_active_vfcmp ? _T_2286 & _T_10 | _T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 &
                _T_4456 : _T_4456;	// sequencer-master.scala:131:52, :183:52
      wire _T_4481 = io_op_bits_active_vfcmp ? _T_2308 & _T_10 | ~_T_10 & _T_4457 : _T_4457;	// sequencer-master.scala:132:52, :184:52
      wire _T_4482 = io_op_bits_active_vfcmp ? _T_2309 & _T_10 | ~_T_10 & _T_4458 : _T_4458;	// sequencer-master.scala:132:52, :184:52
      wire _T_4483 = io_op_bits_active_vfcmp ? _T_2310 & _T_10 | ~_T_10 & _T_4459 : _T_4459;	// sequencer-master.scala:132:52, :184:52
      wire _T_4484 = io_op_bits_active_vfcmp ? _T_2311 & _T_10 | ~_T_10 & _T_4460 : _T_4460;	// sequencer-master.scala:132:52, :184:52
      wire _T_4485 = io_op_bits_active_vfcmp ? _T_2312 & _T_10 | ~_T_10 & _T_4461 : _T_4461;	// sequencer-master.scala:132:52, :184:52
      wire _T_4486 = io_op_bits_active_vfcmp ? _T_2313 & _T_10 | ~_T_10 & _T_4462 : _T_4462;	// sequencer-master.scala:132:52, :184:52
      wire _T_4487 = io_op_bits_active_vfcmp ? _T_2314 & _T_10 | ~_T_10 & _T_4463 : _T_4463;	// sequencer-master.scala:132:52, :184:52
      wire _T_4488 = io_op_bits_active_vfcmp ? _T_2315 & _T_10 | ~_T_10 & _T_4464 : _T_4464;	// sequencer-master.scala:132:52, :184:52
      wire _T_4489 = io_op_bits_active_vfcmp ? _T_2299 & _T_10 | ~_T_10 & _T_4465 : _T_4465;	// sequencer-master.scala:133:52, :185:52
      wire _T_4490 = io_op_bits_active_vfcmp ? _T_2300 & _T_10 | ~_T_10 & _T_4466 : _T_4466;	// sequencer-master.scala:133:52, :185:52
      wire _T_4491 = io_op_bits_active_vfcmp ? _T_2301 & _T_10 | ~_T_10 & _T_4467 : _T_4467;	// sequencer-master.scala:133:52, :185:52
      wire _T_4492 = io_op_bits_active_vfcmp ? _T_2302 & _T_10 | ~_T_10 & _T_4468 : _T_4468;	// sequencer-master.scala:133:52, :185:52
      wire _T_4493 = io_op_bits_active_vfcmp ? _T_2303 & _T_10 | ~_T_10 & _T_4469 : _T_4469;	// sequencer-master.scala:133:52, :185:52
      wire _T_4494 = io_op_bits_active_vfcmp ? _T_2304 & _T_10 | ~_T_10 & _T_4470 : _T_4470;	// sequencer-master.scala:133:52, :185:52
      wire _T_4495 = io_op_bits_active_vfcmp ? _T_2305 & _T_10 | ~_T_10 & _T_4471 : _T_4471;	// sequencer-master.scala:133:52, :185:52
      wire _T_4496 = io_op_bits_active_vfcmp ? _T_2306 & _T_10 | ~_T_10 & _T_4472 : _T_4472;	// sequencer-master.scala:133:52, :185:52
      wire _T_4497 = io_op_bits_active_vfconv ? _T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 & _T_4473 : _T_4473;	// sequencer-master.scala:131:52, :183:52
      wire _T_4498 = io_op_bits_active_vfconv ? _T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 & _T_4474 : _T_4474;	// sequencer-master.scala:131:52, :183:52
      wire _T_4499 = io_op_bits_active_vfconv ? _T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 & _T_4475 : _T_4475;	// sequencer-master.scala:131:52, :183:52
      wire _T_4500 = io_op_bits_active_vfconv ? _T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 & _T_4476 : _T_4476;	// sequencer-master.scala:131:52, :183:52
      wire _T_4501 = io_op_bits_active_vfconv ? _T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 & _T_4477 : _T_4477;	// sequencer-master.scala:131:52, :183:52
      wire _T_4502 = io_op_bits_active_vfconv ? _T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 & _T_4478 : _T_4478;	// sequencer-master.scala:131:52, :183:52
      wire _T_4503 = io_op_bits_active_vfconv ? _T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 & _T_4479 : _T_4479;	// sequencer-master.scala:131:52, :183:52
      wire _T_4504 = io_op_bits_active_vfconv ? _T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 & _T_4480 : _T_4480;	// sequencer-master.scala:131:52, :183:52
      wire _T_4505 = io_op_bits_active_vrpred ? _T_2238 & _T_10 | ~_T_10 & _T_4497 : _T_4497;	// sequencer-master.scala:131:52, :183:52
      wire _T_4506 = io_op_bits_active_vrpred ? _T_2242 & _T_10 | ~_T_10 & _T_4498 : _T_4498;	// sequencer-master.scala:131:52, :183:52
      wire _T_4507 = io_op_bits_active_vrpred ? _T_2246 & _T_10 | ~_T_10 & _T_4499 : _T_4499;	// sequencer-master.scala:131:52, :183:52
      wire _T_4508 = io_op_bits_active_vrpred ? _T_2250 & _T_10 | ~_T_10 & _T_4500 : _T_4500;	// sequencer-master.scala:131:52, :183:52
      wire _T_4509 = io_op_bits_active_vrpred ? _T_2254 & _T_10 | ~_T_10 & _T_4501 : _T_4501;	// sequencer-master.scala:131:52, :183:52
      wire _T_4510 = io_op_bits_active_vrpred ? _T_2258 & _T_10 | ~_T_10 & _T_4502 : _T_4502;	// sequencer-master.scala:131:52, :183:52
      wire _T_4511 = io_op_bits_active_vrpred ? _T_2262 & _T_10 | ~_T_10 & _T_4503 : _T_4503;	// sequencer-master.scala:131:52, :183:52
      wire _T_4512 = io_op_bits_active_vrpred ? _T_2266 & _T_10 | ~_T_10 & _T_4504 : _T_4504;	// sequencer-master.scala:131:52, :183:52
      wire _T_4513 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2308 & _T_10 | ~_T_10 & _T_4481 : _T_4481);	// sequencer-master.scala:132:52, :184:52
      wire _T_4514 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2299 & _T_10 | ~_T_10 & _T_4489 : _T_4489);	// sequencer-master.scala:133:52, :185:52
      wire _T_4515 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2309 & _T_10 | ~_T_10 & _T_4482 : _T_4482);	// sequencer-master.scala:132:52, :184:52
      wire _T_4516 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2300 & _T_10 | ~_T_10 & _T_4490 : _T_4490);	// sequencer-master.scala:133:52, :185:52
      wire _T_4517 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2310 & _T_10 | ~_T_10 & _T_4483 : _T_4483);	// sequencer-master.scala:132:52, :184:52
      wire _T_4518 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2301 & _T_10 | ~_T_10 & _T_4491 : _T_4491);	// sequencer-master.scala:133:52, :185:52
      wire _T_4519 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2311 & _T_10 | ~_T_10 & _T_4484 : _T_4484);	// sequencer-master.scala:132:52, :184:52
      wire _T_4520 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2302 & _T_10 | ~_T_10 & _T_4492 : _T_4492);	// sequencer-master.scala:133:52, :185:52
      wire _T_4521 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2312 & _T_10 | ~_T_10 & _T_4485 : _T_4485);	// sequencer-master.scala:132:52, :184:52
      wire _T_4522 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2303 & _T_10 | ~_T_10 & _T_4493 : _T_4493);	// sequencer-master.scala:133:52, :185:52
      wire _T_4523 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2313 & _T_10 | ~_T_10 & _T_4486 : _T_4486);	// sequencer-master.scala:132:52, :184:52
      wire _T_4524 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2304 & _T_10 | ~_T_10 & _T_4494 : _T_4494);	// sequencer-master.scala:133:52, :185:52
      wire _T_4525 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2314 & _T_10 | ~_T_10 & _T_4487 : _T_4487);	// sequencer-master.scala:132:52, :184:52
      wire _T_4526 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2305 & _T_10 | ~_T_10 & _T_4495 : _T_4495);	// sequencer-master.scala:133:52, :185:52
      wire _T_4527 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2315 & _T_10 | ~_T_10 & _T_4488 : _T_4488);	// sequencer-master.scala:132:52, :184:52
      wire _T_4528 = (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                (io_op_bits_active_vfconv ? _T_2306 & _T_10 | ~_T_10 & _T_4496 : _T_4496);	// sequencer-master.scala:133:52, :185:52
      wire _T_4529 = io_op_bits_active_vrfirst ? _T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 & _T_4505 : _T_4505;	// sequencer-master.scala:131:52, :183:52
      wire _T_4530 = io_op_bits_active_vrfirst ? _T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 & _T_4506 : _T_4506;	// sequencer-master.scala:131:52, :183:52
      wire _T_4531 = io_op_bits_active_vrfirst ? _T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 & _T_4507 : _T_4507;	// sequencer-master.scala:131:52, :183:52
      wire _T_4532 = io_op_bits_active_vrfirst ? _T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 & _T_4508 : _T_4508;	// sequencer-master.scala:131:52, :183:52
      wire _T_4533 = io_op_bits_active_vrfirst ? _T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 & _T_4509 : _T_4509;	// sequencer-master.scala:131:52, :183:52
      wire _T_4534 = io_op_bits_active_vrfirst ? _T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 & _T_4510 : _T_4510;	// sequencer-master.scala:131:52, :183:52
      wire _T_4535 = io_op_bits_active_vrfirst ? _T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 & _T_4511 : _T_4511;	// sequencer-master.scala:131:52, :183:52
      wire _T_4536 = io_op_bits_active_vrfirst ? _T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 & _T_4512 : _T_4512;	// sequencer-master.scala:131:52, :183:52
      wire _T_4537 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_132 | _T_2279 & _T_297 | _T_2238 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2269 & _T_10 | _T_2238 & _T_10 | ~_T_10 & _T_4529)) : _T_4529;	// sequencer-master.scala:131:52, :183:52
      wire _T_4538 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_133 | _T_2280 & _T_297 | _T_2242 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2270 & _T_10 | _T_2242 & _T_10 | ~_T_10 & _T_4530)) : _T_4530;	// sequencer-master.scala:131:52, :183:52
      wire _T_4539 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_134 | _T_2281 & _T_297 | _T_2246 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2271 & _T_10 | _T_2246 & _T_10 | ~_T_10 & _T_4531)) : _T_4531;	// sequencer-master.scala:131:52, :183:52
      wire _T_4540 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_135 | _T_2282 & _T_297 | _T_2250 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2272 & _T_10 | _T_2250 & _T_10 | ~_T_10 & _T_4532)) : _T_4532;	// sequencer-master.scala:131:52, :183:52
      wire _T_4541 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_136 | _T_2283 & _T_297 | _T_2254 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2273 & _T_10 | _T_2254 & _T_10 | ~_T_10 & _T_4533)) : _T_4533;	// sequencer-master.scala:131:52, :183:52
      wire _T_4542 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_137 | _T_2284 & _T_297 | _T_2258 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2274 & _T_10 | _T_2258 & _T_10 | ~_T_10 & _T_4534)) : _T_4534;	// sequencer-master.scala:131:52, :183:52
      wire _T_4543 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & _T_138 | _T_2285 & _T_297 | _T_2262 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2275 & _T_10 | _T_2262 & _T_10 | ~_T_10 & _T_4535)) : _T_4535;	// sequencer-master.scala:131:52, :183:52
      wire _T_4544 = io_op_bits_active_vamo ? ~_T_320 & (_T_297 & &_T_0 | _T_2286 & _T_297 | _T_2266 & _T_297 |
                ~_T_297 & ~_T_138 & (_T_2276 & _T_10 | _T_2266 & _T_10 | ~_T_10 & _T_4536)) : _T_4536;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4545 = io_op_bits_active_vamo ? _T_2308 & _T_320 | ~_T_320 & ~_T_297 & (_T_2308 & _T_138 | ~_T_138
                & ~_T_10 & _T_4513) : _T_4513;	// sequencer-master.scala:132:52, :184:52
      wire _T_4546 = io_op_bits_active_vamo ? _T_2309 & _T_320 | ~_T_320 & ~_T_297 & (_T_2309 & _T_138 | ~_T_138
                & ~_T_10 & _T_4515) : _T_4515;	// sequencer-master.scala:132:52, :184:52
      wire _T_4547 = io_op_bits_active_vamo ? _T_2310 & _T_320 | ~_T_320 & ~_T_297 & (_T_2310 & _T_138 | ~_T_138
                & ~_T_10 & _T_4517) : _T_4517;	// sequencer-master.scala:132:52, :184:52
      wire _T_4548 = io_op_bits_active_vamo ? _T_2311 & _T_320 | ~_T_320 & ~_T_297 & (_T_2311 & _T_138 | ~_T_138
                & ~_T_10 & _T_4519) : _T_4519;	// sequencer-master.scala:132:52, :184:52
      wire _T_4549 = io_op_bits_active_vamo ? _T_2312 & _T_320 | ~_T_320 & ~_T_297 & (_T_2312 & _T_138 | ~_T_138
                & ~_T_10 & _T_4521) : _T_4521;	// sequencer-master.scala:132:52, :184:52
      wire _T_4550 = io_op_bits_active_vamo ? _T_2313 & _T_320 | ~_T_320 & ~_T_297 & (_T_2313 & _T_138 | ~_T_138
                & ~_T_10 & _T_4523) : _T_4523;	// sequencer-master.scala:132:52, :184:52
      wire _T_4551 = io_op_bits_active_vamo ? _T_2314 & _T_320 | ~_T_320 & ~_T_297 & (_T_2314 & _T_138 | ~_T_138
                & ~_T_10 & _T_4525) : _T_4525;	// sequencer-master.scala:132:52, :184:52
      wire _T_4552 = io_op_bits_active_vamo ? _T_2315 & _T_320 | ~_T_320 & ~_T_297 & (_T_2315 & _T_138 | ~_T_138
                & ~_T_10 & _T_4527) : _T_4527;	// sequencer-master.scala:132:52, :184:52
      wire _T_4553 = io_op_bits_active_vamo ? _T_2299 & _T_320 | ~_T_320 & ~_T_297 & (_T_2299 & _T_138 | ~_T_138
                & ~_T_10 & _T_4514) : _T_4514;	// sequencer-master.scala:133:52, :185:52
      wire _T_4554 = io_op_bits_active_vamo ? _T_2300 & _T_320 | ~_T_320 & ~_T_297 & (_T_2300 & _T_138 | ~_T_138
                & ~_T_10 & _T_4516) : _T_4516;	// sequencer-master.scala:133:52, :185:52
      wire _T_4555 = io_op_bits_active_vamo ? _T_2301 & _T_320 | ~_T_320 & ~_T_297 & (_T_2301 & _T_138 | ~_T_138
                & ~_T_10 & _T_4518) : _T_4518;	// sequencer-master.scala:133:52, :185:52
      wire _T_4556 = io_op_bits_active_vamo ? _T_2302 & _T_320 | ~_T_320 & ~_T_297 & (_T_2302 & _T_138 | ~_T_138
                & ~_T_10 & _T_4520) : _T_4520;	// sequencer-master.scala:133:52, :185:52
      wire _T_4557 = io_op_bits_active_vamo ? _T_2303 & _T_320 | ~_T_320 & ~_T_297 & (_T_2303 & _T_138 | ~_T_138
                & ~_T_10 & _T_4522) : _T_4522;	// sequencer-master.scala:133:52, :185:52
      wire _T_4558 = io_op_bits_active_vamo ? _T_2304 & _T_320 | ~_T_320 & ~_T_297 & (_T_2304 & _T_138 | ~_T_138
                & ~_T_10 & _T_4524) : _T_4524;	// sequencer-master.scala:133:52, :185:52
      wire _T_4559 = io_op_bits_active_vamo ? _T_2305 & _T_320 | ~_T_320 & ~_T_297 & (_T_2305 & _T_138 | ~_T_138
                & ~_T_10 & _T_4526) : _T_4526;	// sequencer-master.scala:133:52, :185:52
      wire _T_4560 = io_op_bits_active_vamo ? _T_2306 & _T_320 | ~_T_320 & ~_T_297 & (_T_2306 & _T_138 | ~_T_138
                & ~_T_10 & _T_4528) : _T_4528;	// sequencer-master.scala:133:52, :185:52
      wire _T_4561 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2279 & _T_10 | _T_2238 & _T_10 | ~_T_10 &
                _T_4537) : _T_4537;	// sequencer-master.scala:131:52, :183:52
      wire _T_4562 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2280 & _T_10 | _T_2242 & _T_10 | ~_T_10 &
                _T_4538) : _T_4538;	// sequencer-master.scala:131:52, :183:52
      wire _T_4563 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2281 & _T_10 | _T_2246 & _T_10 | ~_T_10 &
                _T_4539) : _T_4539;	// sequencer-master.scala:131:52, :183:52
      wire _T_4564 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2282 & _T_10 | _T_2250 & _T_10 | ~_T_10 &
                _T_4540) : _T_4540;	// sequencer-master.scala:131:52, :183:52
      wire _T_4565 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2283 & _T_10 | _T_2254 & _T_10 | ~_T_10 &
                _T_4541) : _T_4541;	// sequencer-master.scala:131:52, :183:52
      wire _T_4566 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2284 & _T_10 | _T_2258 & _T_10 | ~_T_10 &
                _T_4542) : _T_4542;	// sequencer-master.scala:131:52, :183:52
      wire _T_4567 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2285 & _T_10 | _T_2262 & _T_10 | ~_T_10 &
                _T_4543) : _T_4543;	// sequencer-master.scala:131:52, :183:52
      wire _T_4568 = io_op_bits_active_vldx ? ~_T_297 & ~_T_138 & (_T_2286 & _T_10 | _T_2266 & _T_10 | ~_T_10 &
                _T_4544) : _T_4544;	// sequencer-master.scala:131:52, :183:52
      wire _T_4569 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2308
                & _T_297 | ~_T_297 & (_T_2308 & _T_138 | ~_T_138 & ~_T_10 & _T_4545) : _T_4545);	// sequencer-master.scala:132:52, :184:52
      wire _T_4570 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2299
                & _T_297 | ~_T_297 & (_T_2299 & _T_138 | ~_T_138 & ~_T_10 & _T_4553) : _T_4553);	// sequencer-master.scala:133:52, :185:52
      wire _T_4571 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2309
                & _T_297 | ~_T_297 & (_T_2309 & _T_138 | ~_T_138 & ~_T_10 & _T_4546) : _T_4546);	// sequencer-master.scala:132:52, :184:52
      wire _T_4572 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2300
                & _T_297 | ~_T_297 & (_T_2300 & _T_138 | ~_T_138 & ~_T_10 & _T_4554) : _T_4554);	// sequencer-master.scala:133:52, :185:52
      wire _T_4573 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2310
                & _T_297 | ~_T_297 & (_T_2310 & _T_138 | ~_T_138 & ~_T_10 & _T_4547) : _T_4547);	// sequencer-master.scala:132:52, :184:52
      wire _T_4574 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2301
                & _T_297 | ~_T_297 & (_T_2301 & _T_138 | ~_T_138 & ~_T_10 & _T_4555) : _T_4555);	// sequencer-master.scala:133:52, :185:52
      wire _T_4575 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2311
                & _T_297 | ~_T_297 & (_T_2311 & _T_138 | ~_T_138 & ~_T_10 & _T_4548) : _T_4548);	// sequencer-master.scala:132:52, :184:52
      wire _T_4576 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2302
                & _T_297 | ~_T_297 & (_T_2302 & _T_138 | ~_T_138 & ~_T_10 & _T_4556) : _T_4556);	// sequencer-master.scala:133:52, :185:52
      wire _T_4577 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2312
                & _T_297 | ~_T_297 & (_T_2312 & _T_138 | ~_T_138 & ~_T_10 & _T_4549) : _T_4549);	// sequencer-master.scala:132:52, :184:52
      wire _T_4578 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2303
                & _T_297 | ~_T_297 & (_T_2303 & _T_138 | ~_T_138 & ~_T_10 & _T_4557) : _T_4557);	// sequencer-master.scala:133:52, :185:52
      wire _T_4579 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2313
                & _T_297 | ~_T_297 & (_T_2313 & _T_138 | ~_T_138 & ~_T_10 & _T_4550) : _T_4550);	// sequencer-master.scala:132:52, :184:52
      wire _T_4580 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2304
                & _T_297 | ~_T_297 & (_T_2304 & _T_138 | ~_T_138 & ~_T_10 & _T_4558) : _T_4558);	// sequencer-master.scala:133:52, :185:52
      wire _T_4581 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2314
                & _T_297 | ~_T_297 & (_T_2314 & _T_138 | ~_T_138 & ~_T_10 & _T_4551) : _T_4551);	// sequencer-master.scala:132:52, :184:52
      wire _T_4582 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2305
                & _T_297 | ~_T_297 & (_T_2305 & _T_138 | ~_T_138 & ~_T_10 & _T_4559) : _T_4559);	// sequencer-master.scala:133:52, :185:52
      wire _T_4583 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2315
                & _T_297 | ~_T_297 & (_T_2315 & _T_138 | ~_T_138 & ~_T_10 & _T_4552) : _T_4552);	// sequencer-master.scala:132:52, :184:52
      wire _T_4584 = (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vldx ? _T_2306
                & _T_297 | ~_T_297 & (_T_2306 & _T_138 | ~_T_138 & ~_T_10 & _T_4560) : _T_4560);	// sequencer-master.scala:133:52, :185:52
      wire _T_4585 = io_op_bits_active_vstx ? _T_297 & _T_132 | _T_2299 & _T_297 | _T_2238 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2279 & _T_10 | _T_2238 & _T_10 | ~_T_10 & _T_4561) : _T_4561;	// sequencer-master.scala:131:52, :183:52
      wire _T_4586 = io_op_bits_active_vstx ? _T_297 & _T_133 | _T_2300 & _T_297 | _T_2242 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2280 & _T_10 | _T_2242 & _T_10 | ~_T_10 & _T_4562) : _T_4562;	// sequencer-master.scala:131:52, :183:52
      wire _T_4587 = io_op_bits_active_vstx ? _T_297 & _T_134 | _T_2301 & _T_297 | _T_2246 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2281 & _T_10 | _T_2246 & _T_10 | ~_T_10 & _T_4563) : _T_4563;	// sequencer-master.scala:131:52, :183:52
      wire _T_4588 = io_op_bits_active_vstx ? _T_297 & _T_135 | _T_2302 & _T_297 | _T_2250 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2282 & _T_10 | _T_2250 & _T_10 | ~_T_10 & _T_4564) : _T_4564;	// sequencer-master.scala:131:52, :183:52
      wire _T_4589 = io_op_bits_active_vstx ? _T_297 & _T_136 | _T_2303 & _T_297 | _T_2254 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2283 & _T_10 | _T_2254 & _T_10 | ~_T_10 & _T_4565) : _T_4565;	// sequencer-master.scala:131:52, :183:52
      wire _T_4590 = io_op_bits_active_vstx ? _T_297 & _T_137 | _T_2304 & _T_297 | _T_2258 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2284 & _T_10 | _T_2258 & _T_10 | ~_T_10 & _T_4566) : _T_4566;	// sequencer-master.scala:131:52, :183:52
      wire _T_4591 = io_op_bits_active_vstx ? _T_297 & _T_138 | _T_2305 & _T_297 | _T_2262 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2285 & _T_10 | _T_2262 & _T_10 | ~_T_10 & _T_4567) : _T_4567;	// sequencer-master.scala:131:52, :183:52
      wire _T_4592 = io_op_bits_active_vstx ? _T_297 & &_T_0 | _T_2306 & _T_297 | _T_2266 & _T_297 | ~_T_297 &
                ~_T_138 & (_T_2286 & _T_10 | _T_2266 & _T_10 | ~_T_10 & _T_4568) : _T_4568;	// sequencer-master.scala:131:52, :183:52, :267:35
      wire _T_4593 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2238 & _T_10 | ~_T_10 & _T_4585) : _T_4585;	// sequencer-master.scala:131:52, :183:52
      wire _T_4594 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2242 & _T_10 | ~_T_10 & _T_4586) : _T_4586;	// sequencer-master.scala:131:52, :183:52
      wire _T_4595 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2246 & _T_10 | ~_T_10 & _T_4587) : _T_4587;	// sequencer-master.scala:131:52, :183:52
      wire _T_4596 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2250 & _T_10 | ~_T_10 & _T_4588) : _T_4588;	// sequencer-master.scala:131:52, :183:52
      wire _T_4597 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2254 & _T_10 | ~_T_10 & _T_4589) : _T_4589;	// sequencer-master.scala:131:52, :183:52
      wire _T_4598 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2258 & _T_10 | ~_T_10 & _T_4590) : _T_4590;	// sequencer-master.scala:131:52, :183:52
      wire _T_4599 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2262 & _T_10 | ~_T_10 & _T_4591) : _T_4591;	// sequencer-master.scala:131:52, :183:52
      wire _T_4600 = io_op_bits_active_vld ? ~_T_297 & ~_T_138 & (_T_2266 & _T_10 | ~_T_10 & _T_4592) : _T_4592;	// sequencer-master.scala:131:52, :183:52
      wire _T_4601 = io_op_bits_active_vint ? _T_2279 & &tail | _T_2269 & &tail | _T_2238 & &tail | ~(&tail) &
                e_7_raw_0 : e_7_raw_0;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4602 = io_op_bits_active_vint ? _T_2280 & &tail | _T_2270 & &tail | _T_2242 & &tail | ~(&tail) &
                e_7_raw_1 : e_7_raw_1;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4603 = io_op_bits_active_vint ? _T_2281 & &tail | _T_2271 & &tail | _T_2246 & &tail | ~(&tail) &
                e_7_raw_2 : e_7_raw_2;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4604 = io_op_bits_active_vint ? _T_2282 & &tail | _T_2272 & &tail | _T_2250 & &tail | ~(&tail) &
                e_7_raw_3 : e_7_raw_3;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4605 = io_op_bits_active_vint ? _T_2283 & &tail | _T_2273 & &tail | _T_2254 & &tail | ~(&tail) &
                e_7_raw_4 : e_7_raw_4;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4606 = io_op_bits_active_vint ? _T_2284 & &tail | _T_2274 & &tail | _T_2258 & &tail | ~(&tail) &
                e_7_raw_5 : e_7_raw_5;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4607 = io_op_bits_active_vint ? _T_2285 & &tail | _T_2275 & &tail | _T_2262 & &tail | ~(&tail) &
                e_7_raw_6 : e_7_raw_6;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4608 = io_op_bits_active_vint ? _T_2286 & &tail | _T_2276 & &tail | _T_2266 & &tail | ~(&tail) &
                e_7_raw_7 : e_7_raw_7;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4609 = io_op_bits_active_vint ? _T_2308 & &tail | ~(&tail) & e_7_war_0 : e_7_war_0;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4610 = io_op_bits_active_vint ? _T_2309 & &tail | ~(&tail) & e_7_war_1 : e_7_war_1;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4611 = io_op_bits_active_vint ? _T_2310 & &tail | ~(&tail) & e_7_war_2 : e_7_war_2;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4612 = io_op_bits_active_vint ? _T_2311 & &tail | ~(&tail) & e_7_war_3 : e_7_war_3;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4613 = io_op_bits_active_vint ? _T_2312 & &tail | ~(&tail) & e_7_war_4 : e_7_war_4;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4614 = io_op_bits_active_vint ? _T_2313 & &tail | ~(&tail) & e_7_war_5 : e_7_war_5;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4615 = io_op_bits_active_vint ? _T_2314 & &tail | ~(&tail) & e_7_war_6 : e_7_war_6;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4616 = io_op_bits_active_vint ? _T_2315 & &tail | ~(&tail) & e_7_war_7 : e_7_war_7;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4617 = io_op_bits_active_vint ? _T_2299 & &tail | ~(&tail) & e_7_waw_0 : e_7_waw_0;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4618 = io_op_bits_active_vint ? _T_2300 & &tail | ~(&tail) & e_7_waw_1 : e_7_waw_1;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4619 = io_op_bits_active_vint ? _T_2301 & &tail | ~(&tail) & e_7_waw_2 : e_7_waw_2;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4620 = io_op_bits_active_vint ? _T_2302 & &tail | ~(&tail) & e_7_waw_3 : e_7_waw_3;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4621 = io_op_bits_active_vint ? _T_2303 & &tail | ~(&tail) & e_7_waw_4 : e_7_waw_4;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4622 = io_op_bits_active_vint ? _T_2304 & &tail | ~(&tail) & e_7_waw_5 : e_7_waw_5;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4623 = io_op_bits_active_vint ? _T_2305 & &tail | ~(&tail) & e_7_waw_6 : e_7_waw_6;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4624 = io_op_bits_active_vint ? _T_2306 & &tail | ~(&tail) & e_7_waw_7 : e_7_waw_7;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4625 = io_op_bits_active_vipred ? _T_2289 & &tail | _T_2279 & &tail | _T_2269 & &tail | ~(&tail) &
                _T_4601 : _T_4601;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4626 = io_op_bits_active_vipred ? _T_2290 & &tail | _T_2280 & &tail | _T_2270 & &tail | ~(&tail) &
                _T_4602 : _T_4602;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4627 = io_op_bits_active_vipred ? _T_2291 & &tail | _T_2281 & &tail | _T_2271 & &tail | ~(&tail) &
                _T_4603 : _T_4603;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4628 = io_op_bits_active_vipred ? _T_2292 & &tail | _T_2282 & &tail | _T_2272 & &tail | ~(&tail) &
                _T_4604 : _T_4604;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4629 = io_op_bits_active_vipred ? _T_2293 & &tail | _T_2283 & &tail | _T_2273 & &tail | ~(&tail) &
                _T_4605 : _T_4605;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4630 = io_op_bits_active_vipred ? _T_2294 & &tail | _T_2284 & &tail | _T_2274 & &tail | ~(&tail) &
                _T_4606 : _T_4606;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4631 = io_op_bits_active_vipred ? _T_2295 & &tail | _T_2285 & &tail | _T_2275 & &tail | ~(&tail) &
                _T_4607 : _T_4607;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4632 = io_op_bits_active_vipred ? _T_2296 & &tail | _T_2286 & &tail | _T_2276 & &tail | ~(&tail) &
                _T_4608 : _T_4608;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4633 = io_op_bits_active_vipred ? _T_2308 & &tail | ~(&tail) & _T_4609 : _T_4609;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4634 = io_op_bits_active_vipred ? _T_2309 & &tail | ~(&tail) & _T_4610 : _T_4610;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4635 = io_op_bits_active_vipred ? _T_2310 & &tail | ~(&tail) & _T_4611 : _T_4611;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4636 = io_op_bits_active_vipred ? _T_2311 & &tail | ~(&tail) & _T_4612 : _T_4612;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4637 = io_op_bits_active_vipred ? _T_2312 & &tail | ~(&tail) & _T_4613 : _T_4613;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4638 = io_op_bits_active_vipred ? _T_2313 & &tail | ~(&tail) & _T_4614 : _T_4614;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4639 = io_op_bits_active_vipred ? _T_2314 & &tail | ~(&tail) & _T_4615 : _T_4615;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4640 = io_op_bits_active_vipred ? _T_2315 & &tail | ~(&tail) & _T_4616 : _T_4616;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4641 = io_op_bits_active_vipred ? _T_2299 & &tail | ~(&tail) & _T_4617 : _T_4617;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4642 = io_op_bits_active_vipred ? _T_2300 & &tail | ~(&tail) & _T_4618 : _T_4618;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4643 = io_op_bits_active_vipred ? _T_2301 & &tail | ~(&tail) & _T_4619 : _T_4619;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4644 = io_op_bits_active_vipred ? _T_2302 & &tail | ~(&tail) & _T_4620 : _T_4620;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4645 = io_op_bits_active_vipred ? _T_2303 & &tail | ~(&tail) & _T_4621 : _T_4621;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4646 = io_op_bits_active_vipred ? _T_2304 & &tail | ~(&tail) & _T_4622 : _T_4622;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4647 = io_op_bits_active_vipred ? _T_2305 & &tail | ~(&tail) & _T_4623 : _T_4623;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4648 = io_op_bits_active_vipred ? _T_2306 & &tail | ~(&tail) & _T_4624 : _T_4624;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4649 = io_op_bits_active_vimul ? _T_2279 & &tail | _T_2269 & &tail | _T_2238 & &tail | ~(&tail) &
                _T_4625 : _T_4625;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4650 = io_op_bits_active_vimul ? _T_2280 & &tail | _T_2270 & &tail | _T_2242 & &tail | ~(&tail) &
                _T_4626 : _T_4626;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4651 = io_op_bits_active_vimul ? _T_2281 & &tail | _T_2271 & &tail | _T_2246 & &tail | ~(&tail) &
                _T_4627 : _T_4627;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4652 = io_op_bits_active_vimul ? _T_2282 & &tail | _T_2272 & &tail | _T_2250 & &tail | ~(&tail) &
                _T_4628 : _T_4628;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4653 = io_op_bits_active_vimul ? _T_2283 & &tail | _T_2273 & &tail | _T_2254 & &tail | ~(&tail) &
                _T_4629 : _T_4629;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4654 = io_op_bits_active_vimul ? _T_2284 & &tail | _T_2274 & &tail | _T_2258 & &tail | ~(&tail) &
                _T_4630 : _T_4630;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4655 = io_op_bits_active_vimul ? _T_2285 & &tail | _T_2275 & &tail | _T_2262 & &tail | ~(&tail) &
                _T_4631 : _T_4631;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4656 = io_op_bits_active_vimul ? _T_2286 & &tail | _T_2276 & &tail | _T_2266 & &tail | ~(&tail) &
                _T_4632 : _T_4632;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4657 = io_op_bits_active_vimul ? _T_2308 & &tail | ~(&tail) & _T_4633 : _T_4633;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4658 = io_op_bits_active_vimul ? _T_2309 & &tail | ~(&tail) & _T_4634 : _T_4634;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4659 = io_op_bits_active_vimul ? _T_2310 & &tail | ~(&tail) & _T_4635 : _T_4635;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4660 = io_op_bits_active_vimul ? _T_2311 & &tail | ~(&tail) & _T_4636 : _T_4636;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4661 = io_op_bits_active_vimul ? _T_2312 & &tail | ~(&tail) & _T_4637 : _T_4637;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4662 = io_op_bits_active_vimul ? _T_2313 & &tail | ~(&tail) & _T_4638 : _T_4638;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4663 = io_op_bits_active_vimul ? _T_2314 & &tail | ~(&tail) & _T_4639 : _T_4639;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4664 = io_op_bits_active_vimul ? _T_2315 & &tail | ~(&tail) & _T_4640 : _T_4640;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4665 = io_op_bits_active_vimul ? _T_2299 & &tail | ~(&tail) & _T_4641 : _T_4641;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4666 = io_op_bits_active_vimul ? _T_2300 & &tail | ~(&tail) & _T_4642 : _T_4642;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4667 = io_op_bits_active_vimul ? _T_2301 & &tail | ~(&tail) & _T_4643 : _T_4643;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4668 = io_op_bits_active_vimul ? _T_2302 & &tail | ~(&tail) & _T_4644 : _T_4644;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4669 = io_op_bits_active_vimul ? _T_2303 & &tail | ~(&tail) & _T_4645 : _T_4645;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4670 = io_op_bits_active_vimul ? _T_2304 & &tail | ~(&tail) & _T_4646 : _T_4646;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4671 = io_op_bits_active_vimul ? _T_2305 & &tail | ~(&tail) & _T_4647 : _T_4647;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4672 = io_op_bits_active_vimul ? _T_2306 & &tail | ~(&tail) & _T_4648 : _T_4648;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4673 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2279 & &tail | _T_2269 & &tail | _T_2238 & &tail |
                ~(&tail) & _T_4649) : _T_4649;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4674 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2280 & &tail | _T_2270 & &tail | _T_2242 & &tail |
                ~(&tail) & _T_4650) : _T_4650;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4675 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2281 & &tail | _T_2271 & &tail | _T_2246 & &tail |
                ~(&tail) & _T_4651) : _T_4651;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4676 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2282 & &tail | _T_2272 & &tail | _T_2250 & &tail |
                ~(&tail) & _T_4652) : _T_4652;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4677 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2283 & &tail | _T_2273 & &tail | _T_2254 & &tail |
                ~(&tail) & _T_4653) : _T_4653;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4678 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2284 & &tail | _T_2274 & &tail | _T_2258 & &tail |
                ~(&tail) & _T_4654) : _T_4654;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4679 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2285 & &tail | _T_2275 & &tail | _T_2262 & &tail |
                ~(&tail) & _T_4655) : _T_4655;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4680 = io_op_bits_active_vidiv ? ~(&_T_0) & (_T_2286 & &tail | _T_2276 & &tail | _T_2266 & &tail |
                ~(&tail) & _T_4656) : _T_4656;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4681 = io_op_bits_active_vidiv ? _T_2308 & &_T_0 | ~(&_T_0) & (_T_2308 & &tail | ~(&tail) &
                _T_4657) : _T_4657;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4682 = io_op_bits_active_vidiv ? _T_2309 & &_T_0 | ~(&_T_0) & (_T_2309 & &tail | ~(&tail) &
                _T_4658) : _T_4658;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4683 = io_op_bits_active_vidiv ? _T_2310 & &_T_0 | ~(&_T_0) & (_T_2310 & &tail | ~(&tail) &
                _T_4659) : _T_4659;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4684 = io_op_bits_active_vidiv ? _T_2311 & &_T_0 | ~(&_T_0) & (_T_2311 & &tail | ~(&tail) &
                _T_4660) : _T_4660;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4685 = io_op_bits_active_vidiv ? _T_2312 & &_T_0 | ~(&_T_0) & (_T_2312 & &tail | ~(&tail) &
                _T_4661) : _T_4661;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4686 = io_op_bits_active_vidiv ? _T_2313 & &_T_0 | ~(&_T_0) & (_T_2313 & &tail | ~(&tail) &
                _T_4662) : _T_4662;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4687 = io_op_bits_active_vidiv ? _T_2314 & &_T_0 | ~(&_T_0) & (_T_2314 & &tail | ~(&tail) &
                _T_4663) : _T_4663;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4688 = io_op_bits_active_vidiv ? _T_2315 & &_T_0 | ~(&_T_0) & (_T_2315 & &tail | ~(&tail) &
                _T_4664) : _T_4664;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4689 = io_op_bits_active_vidiv ? _T_2299 & &_T_0 | ~(&_T_0) & (_T_2299 & &tail | ~(&tail) &
                _T_4665) : _T_4665;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4690 = io_op_bits_active_vidiv ? _T_2300 & &_T_0 | ~(&_T_0) & (_T_2300 & &tail | ~(&tail) &
                _T_4666) : _T_4666;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4691 = io_op_bits_active_vidiv ? _T_2301 & &_T_0 | ~(&_T_0) & (_T_2301 & &tail | ~(&tail) &
                _T_4667) : _T_4667;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4692 = io_op_bits_active_vidiv ? _T_2302 & &_T_0 | ~(&_T_0) & (_T_2302 & &tail | ~(&tail) &
                _T_4668) : _T_4668;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4693 = io_op_bits_active_vidiv ? _T_2303 & &_T_0 | ~(&_T_0) & (_T_2303 & &tail | ~(&tail) &
                _T_4669) : _T_4669;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4694 = io_op_bits_active_vidiv ? _T_2304 & &_T_0 | ~(&_T_0) & (_T_2304 & &tail | ~(&tail) &
                _T_4670) : _T_4670;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4695 = io_op_bits_active_vidiv ? _T_2305 & &_T_0 | ~(&_T_0) & (_T_2305 & &tail | ~(&tail) &
                _T_4671) : _T_4671;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4696 = io_op_bits_active_vidiv ? _T_2306 & &_T_0 | ~(&_T_0) & (_T_2306 & &tail | ~(&tail) &
                _T_4672) : _T_4672;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4697 = io_op_bits_active_vfma ? _T_2289 & &tail | _T_2279 & &tail | _T_2269 & &tail | _T_2238 &
                &tail | ~(&tail) & _T_4673 : _T_4673;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4698 = io_op_bits_active_vfma ? _T_2290 & &tail | _T_2280 & &tail | _T_2270 & &tail | _T_2242 &
                &tail | ~(&tail) & _T_4674 : _T_4674;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4699 = io_op_bits_active_vfma ? _T_2291 & &tail | _T_2281 & &tail | _T_2271 & &tail | _T_2246 &
                &tail | ~(&tail) & _T_4675 : _T_4675;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4700 = io_op_bits_active_vfma ? _T_2292 & &tail | _T_2282 & &tail | _T_2272 & &tail | _T_2250 &
                &tail | ~(&tail) & _T_4676 : _T_4676;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4701 = io_op_bits_active_vfma ? _T_2293 & &tail | _T_2283 & &tail | _T_2273 & &tail | _T_2254 &
                &tail | ~(&tail) & _T_4677 : _T_4677;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4702 = io_op_bits_active_vfma ? _T_2294 & &tail | _T_2284 & &tail | _T_2274 & &tail | _T_2258 &
                &tail | ~(&tail) & _T_4678 : _T_4678;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4703 = io_op_bits_active_vfma ? _T_2295 & &tail | _T_2285 & &tail | _T_2275 & &tail | _T_2262 &
                &tail | ~(&tail) & _T_4679 : _T_4679;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4704 = io_op_bits_active_vfma ? _T_2296 & &tail | _T_2286 & &tail | _T_2276 & &tail | _T_2266 &
                &tail | ~(&tail) & _T_4680 : _T_4680;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4705 = io_op_bits_active_vfma ? _T_2308 & &tail | ~(&tail) & _T_4681 : _T_4681;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4706 = io_op_bits_active_vfma ? _T_2309 & &tail | ~(&tail) & _T_4682 : _T_4682;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4707 = io_op_bits_active_vfma ? _T_2310 & &tail | ~(&tail) & _T_4683 : _T_4683;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4708 = io_op_bits_active_vfma ? _T_2311 & &tail | ~(&tail) & _T_4684 : _T_4684;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4709 = io_op_bits_active_vfma ? _T_2312 & &tail | ~(&tail) & _T_4685 : _T_4685;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4710 = io_op_bits_active_vfma ? _T_2313 & &tail | ~(&tail) & _T_4686 : _T_4686;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4711 = io_op_bits_active_vfma ? _T_2314 & &tail | ~(&tail) & _T_4687 : _T_4687;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4712 = io_op_bits_active_vfma ? _T_2315 & &tail | ~(&tail) & _T_4688 : _T_4688;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4713 = io_op_bits_active_vfma ? _T_2299 & &tail | ~(&tail) & _T_4689 : _T_4689;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4714 = io_op_bits_active_vfma ? _T_2300 & &tail | ~(&tail) & _T_4690 : _T_4690;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4715 = io_op_bits_active_vfma ? _T_2301 & &tail | ~(&tail) & _T_4691 : _T_4691;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4716 = io_op_bits_active_vfma ? _T_2302 & &tail | ~(&tail) & _T_4692 : _T_4692;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4717 = io_op_bits_active_vfma ? _T_2303 & &tail | ~(&tail) & _T_4693 : _T_4693;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4718 = io_op_bits_active_vfma ? _T_2304 & &tail | ~(&tail) & _T_4694 : _T_4694;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4719 = io_op_bits_active_vfma ? _T_2305 & &tail | ~(&tail) & _T_4695 : _T_4695;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4720 = io_op_bits_active_vfma ? _T_2306 & &tail | ~(&tail) & _T_4696 : _T_4696;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4721 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2279 & &tail | _T_2269 & &tail | _T_2238 & &tail |
                ~(&tail) & _T_4697) : _T_4697;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4722 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2280 & &tail | _T_2270 & &tail | _T_2242 & &tail |
                ~(&tail) & _T_4698) : _T_4698;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4723 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2281 & &tail | _T_2271 & &tail | _T_2246 & &tail |
                ~(&tail) & _T_4699) : _T_4699;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4724 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2282 & &tail | _T_2272 & &tail | _T_2250 & &tail |
                ~(&tail) & _T_4700) : _T_4700;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4725 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2283 & &tail | _T_2273 & &tail | _T_2254 & &tail |
                ~(&tail) & _T_4701) : _T_4701;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4726 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2284 & &tail | _T_2274 & &tail | _T_2258 & &tail |
                ~(&tail) & _T_4702) : _T_4702;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4727 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2285 & &tail | _T_2275 & &tail | _T_2262 & &tail |
                ~(&tail) & _T_4703) : _T_4703;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4728 = io_op_bits_active_vfdiv ? ~(&_T_0) & (_T_2286 & &tail | _T_2276 & &tail | _T_2266 & &tail |
                ~(&tail) & _T_4704) : _T_4704;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4729 = io_op_bits_active_vfdiv ? _T_2308 & &_T_0 | ~(&_T_0) & (_T_2308 & &tail | ~(&tail) &
                _T_4705) : _T_4705;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4730 = io_op_bits_active_vfdiv ? _T_2309 & &_T_0 | ~(&_T_0) & (_T_2309 & &tail | ~(&tail) &
                _T_4706) : _T_4706;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4731 = io_op_bits_active_vfdiv ? _T_2310 & &_T_0 | ~(&_T_0) & (_T_2310 & &tail | ~(&tail) &
                _T_4707) : _T_4707;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4732 = io_op_bits_active_vfdiv ? _T_2311 & &_T_0 | ~(&_T_0) & (_T_2311 & &tail | ~(&tail) &
                _T_4708) : _T_4708;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4733 = io_op_bits_active_vfdiv ? _T_2312 & &_T_0 | ~(&_T_0) & (_T_2312 & &tail | ~(&tail) &
                _T_4709) : _T_4709;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4734 = io_op_bits_active_vfdiv ? _T_2313 & &_T_0 | ~(&_T_0) & (_T_2313 & &tail | ~(&tail) &
                _T_4710) : _T_4710;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4735 = io_op_bits_active_vfdiv ? _T_2314 & &_T_0 | ~(&_T_0) & (_T_2314 & &tail | ~(&tail) &
                _T_4711) : _T_4711;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4736 = io_op_bits_active_vfdiv ? _T_2315 & &_T_0 | ~(&_T_0) & (_T_2315 & &tail | ~(&tail) &
                _T_4712) : _T_4712;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4737 = io_op_bits_active_vfdiv ? _T_2299 & &_T_0 | ~(&_T_0) & (_T_2299 & &tail | ~(&tail) &
                _T_4713) : _T_4713;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4738 = io_op_bits_active_vfdiv ? _T_2300 & &_T_0 | ~(&_T_0) & (_T_2300 & &tail | ~(&tail) &
                _T_4714) : _T_4714;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4739 = io_op_bits_active_vfdiv ? _T_2301 & &_T_0 | ~(&_T_0) & (_T_2301 & &tail | ~(&tail) &
                _T_4715) : _T_4715;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4740 = io_op_bits_active_vfdiv ? _T_2302 & &_T_0 | ~(&_T_0) & (_T_2302 & &tail | ~(&tail) &
                _T_4716) : _T_4716;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4741 = io_op_bits_active_vfdiv ? _T_2303 & &_T_0 | ~(&_T_0) & (_T_2303 & &tail | ~(&tail) &
                _T_4717) : _T_4717;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4742 = io_op_bits_active_vfdiv ? _T_2304 & &_T_0 | ~(&_T_0) & (_T_2304 & &tail | ~(&tail) &
                _T_4718) : _T_4718;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4743 = io_op_bits_active_vfdiv ? _T_2305 & &_T_0 | ~(&_T_0) & (_T_2305 & &tail | ~(&tail) &
                _T_4719) : _T_4719;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4744 = io_op_bits_active_vfdiv ? _T_2306 & &_T_0 | ~(&_T_0) & (_T_2306 & &tail | ~(&tail) &
                _T_4720) : _T_4720;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4745 = io_op_bits_active_vfcmp ? _T_2279 & &tail | _T_2269 & &tail | _T_2238 & &tail | ~(&tail) &
                _T_4721 : _T_4721;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4746 = io_op_bits_active_vfcmp ? _T_2280 & &tail | _T_2270 & &tail | _T_2242 & &tail | ~(&tail) &
                _T_4722 : _T_4722;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4747 = io_op_bits_active_vfcmp ? _T_2281 & &tail | _T_2271 & &tail | _T_2246 & &tail | ~(&tail) &
                _T_4723 : _T_4723;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4748 = io_op_bits_active_vfcmp ? _T_2282 & &tail | _T_2272 & &tail | _T_2250 & &tail | ~(&tail) &
                _T_4724 : _T_4724;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4749 = io_op_bits_active_vfcmp ? _T_2283 & &tail | _T_2273 & &tail | _T_2254 & &tail | ~(&tail) &
                _T_4725 : _T_4725;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4750 = io_op_bits_active_vfcmp ? _T_2284 & &tail | _T_2274 & &tail | _T_2258 & &tail | ~(&tail) &
                _T_4726 : _T_4726;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4751 = io_op_bits_active_vfcmp ? _T_2285 & &tail | _T_2275 & &tail | _T_2262 & &tail | ~(&tail) &
                _T_4727 : _T_4727;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4752 = io_op_bits_active_vfcmp ? _T_2286 & &tail | _T_2276 & &tail | _T_2266 & &tail | ~(&tail) &
                _T_4728 : _T_4728;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4753 = io_op_bits_active_vfcmp ? _T_2308 & &tail | ~(&tail) & _T_4729 : _T_4729;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4754 = io_op_bits_active_vfcmp ? _T_2309 & &tail | ~(&tail) & _T_4730 : _T_4730;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4755 = io_op_bits_active_vfcmp ? _T_2310 & &tail | ~(&tail) & _T_4731 : _T_4731;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4756 = io_op_bits_active_vfcmp ? _T_2311 & &tail | ~(&tail) & _T_4732 : _T_4732;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4757 = io_op_bits_active_vfcmp ? _T_2312 & &tail | ~(&tail) & _T_4733 : _T_4733;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4758 = io_op_bits_active_vfcmp ? _T_2313 & &tail | ~(&tail) & _T_4734 : _T_4734;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4759 = io_op_bits_active_vfcmp ? _T_2314 & &tail | ~(&tail) & _T_4735 : _T_4735;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4760 = io_op_bits_active_vfcmp ? _T_2315 & &tail | ~(&tail) & _T_4736 : _T_4736;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4761 = io_op_bits_active_vfcmp ? _T_2299 & &tail | ~(&tail) & _T_4737 : _T_4737;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4762 = io_op_bits_active_vfcmp ? _T_2300 & &tail | ~(&tail) & _T_4738 : _T_4738;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4763 = io_op_bits_active_vfcmp ? _T_2301 & &tail | ~(&tail) & _T_4739 : _T_4739;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4764 = io_op_bits_active_vfcmp ? _T_2302 & &tail | ~(&tail) & _T_4740 : _T_4740;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4765 = io_op_bits_active_vfcmp ? _T_2303 & &tail | ~(&tail) & _T_4741 : _T_4741;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4766 = io_op_bits_active_vfcmp ? _T_2304 & &tail | ~(&tail) & _T_4742 : _T_4742;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4767 = io_op_bits_active_vfcmp ? _T_2305 & &tail | ~(&tail) & _T_4743 : _T_4743;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4768 = io_op_bits_active_vfcmp ? _T_2306 & &tail | ~(&tail) & _T_4744 : _T_4744;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4769 = io_op_bits_active_vfconv ? _T_2269 & &tail | _T_2238 & &tail | ~(&tail) & _T_4745 : _T_4745;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4770 = io_op_bits_active_vfconv ? _T_2270 & &tail | _T_2242 & &tail | ~(&tail) & _T_4746 : _T_4746;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4771 = io_op_bits_active_vfconv ? _T_2271 & &tail | _T_2246 & &tail | ~(&tail) & _T_4747 : _T_4747;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4772 = io_op_bits_active_vfconv ? _T_2272 & &tail | _T_2250 & &tail | ~(&tail) & _T_4748 : _T_4748;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4773 = io_op_bits_active_vfconv ? _T_2273 & &tail | _T_2254 & &tail | ~(&tail) & _T_4749 : _T_4749;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4774 = io_op_bits_active_vfconv ? _T_2274 & &tail | _T_2258 & &tail | ~(&tail) & _T_4750 : _T_4750;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4775 = io_op_bits_active_vfconv ? _T_2275 & &tail | _T_2262 & &tail | ~(&tail) & _T_4751 : _T_4751;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4776 = io_op_bits_active_vfconv ? _T_2276 & &tail | _T_2266 & &tail | ~(&tail) & _T_4752 : _T_4752;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4777 = io_op_bits_active_vrpred ? _T_2238 & &tail | ~(&tail) & _T_4769 : _T_4769;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4778 = io_op_bits_active_vrpred ? _T_2242 & &tail | ~(&tail) & _T_4770 : _T_4770;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4779 = io_op_bits_active_vrpred ? _T_2246 & &tail | ~(&tail) & _T_4771 : _T_4771;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4780 = io_op_bits_active_vrpred ? _T_2250 & &tail | ~(&tail) & _T_4772 : _T_4772;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4781 = io_op_bits_active_vrpred ? _T_2254 & &tail | ~(&tail) & _T_4773 : _T_4773;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4782 = io_op_bits_active_vrpred ? _T_2258 & &tail | ~(&tail) & _T_4774 : _T_4774;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4783 = io_op_bits_active_vrpred ? _T_2262 & &tail | ~(&tail) & _T_4775 : _T_4775;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4784 = io_op_bits_active_vrpred ? _T_2266 & &tail | ~(&tail) & _T_4776 : _T_4776;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4785 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2308 & &tail | ~(&tail) & _T_4753 : _T_4753);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4786 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2299 & &tail | ~(&tail) & _T_4761 : _T_4761);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4787 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2309 & &tail | ~(&tail) & _T_4754 : _T_4754);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4788 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2300 & &tail | ~(&tail) & _T_4762 : _T_4762);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4789 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2310 & &tail | ~(&tail) & _T_4755 : _T_4755);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4790 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2301 & &tail | ~(&tail) & _T_4763 : _T_4763);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4791 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2311 & &tail | ~(&tail) & _T_4756 : _T_4756);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4792 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2302 & &tail | ~(&tail) & _T_4764 : _T_4764);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4793 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2312 & &tail | ~(&tail) & _T_4757 : _T_4757);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4794 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2303 & &tail | ~(&tail) & _T_4765 : _T_4765);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4795 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2313 & &tail | ~(&tail) & _T_4758 : _T_4758);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4796 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2304 & &tail | ~(&tail) & _T_4766 : _T_4766);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4797 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2314 & &tail | ~(&tail) & _T_4759 : _T_4759);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4798 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2305 & &tail | ~(&tail) & _T_4767 : _T_4767);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4799 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2315 & &tail | ~(&tail) & _T_4760 : _T_4760);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4800 = (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                (io_op_bits_active_vfconv ? _T_2306 & &tail | ~(&tail) & _T_4768 : _T_4768);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4801 = io_op_bits_active_vrfirst ? _T_2269 & &tail | _T_2238 & &tail | ~(&tail) & _T_4777 :
                _T_4777;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4802 = io_op_bits_active_vrfirst ? _T_2270 & &tail | _T_2242 & &tail | ~(&tail) & _T_4778 :
                _T_4778;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4803 = io_op_bits_active_vrfirst ? _T_2271 & &tail | _T_2246 & &tail | ~(&tail) & _T_4779 :
                _T_4779;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4804 = io_op_bits_active_vrfirst ? _T_2272 & &tail | _T_2250 & &tail | ~(&tail) & _T_4780 :
                _T_4780;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4805 = io_op_bits_active_vrfirst ? _T_2273 & &tail | _T_2254 & &tail | ~(&tail) & _T_4781 :
                _T_4781;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4806 = io_op_bits_active_vrfirst ? _T_2274 & &tail | _T_2258 & &tail | ~(&tail) & _T_4782 :
                _T_4782;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4807 = io_op_bits_active_vrfirst ? _T_2275 & &tail | _T_2262 & &tail | ~(&tail) & _T_4783 :
                _T_4783;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4808 = io_op_bits_active_vrfirst ? _T_2276 & &tail | _T_2266 & &tail | ~(&tail) & _T_4784 :
                _T_4784;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4809 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_132 | _T_2279 & &_T_1 | _T_2238 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2269 & &tail | _T_2238 & &tail | ~(&tail) & _T_4801)) : _T_4801;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4810 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_133 | _T_2280 & &_T_1 | _T_2242 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2270 & &tail | _T_2242 & &tail | ~(&tail) & _T_4802)) : _T_4802;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4811 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_134 | _T_2281 & &_T_1 | _T_2246 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2271 & &tail | _T_2246 & &tail | ~(&tail) & _T_4803)) : _T_4803;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4812 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_135 | _T_2282 & &_T_1 | _T_2250 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2272 & &tail | _T_2250 & &tail | ~(&tail) & _T_4804)) : _T_4804;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4813 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_136 | _T_2283 & &_T_1 | _T_2254 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2273 & &tail | _T_2254 & &tail | ~(&tail) & _T_4805)) : _T_4805;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4814 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_137 | _T_2284 & &_T_1 | _T_2258 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2274 & &tail | _T_2258 & &tail | ~(&tail) & _T_4806)) : _T_4806;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4815 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & _T_138 | _T_2285 & &_T_1 | _T_2262 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2275 & &tail | _T_2262 & &tail | ~(&tail) & _T_4807)) : _T_4807;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4816 = io_op_bits_active_vamo ? ~(&_T_2) & (&_T_1 & &_T_0 | _T_2286 & &_T_1 | _T_2266 & &_T_1 |
                ~(&_T_1) & ~(&_T_0) & (_T_2276 & &tail | _T_2266 & &tail | ~(&tail) & _T_4808)) : _T_4808;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4817 = io_op_bits_active_vamo ? _T_2308 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2308 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4785) : _T_4785;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4818 = io_op_bits_active_vamo ? _T_2309 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2309 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4787) : _T_4787;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4819 = io_op_bits_active_vamo ? _T_2310 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2310 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4789) : _T_4789;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4820 = io_op_bits_active_vamo ? _T_2311 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2311 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4791) : _T_4791;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4821 = io_op_bits_active_vamo ? _T_2312 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2312 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4793) : _T_4793;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4822 = io_op_bits_active_vamo ? _T_2313 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2313 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4795) : _T_4795;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4823 = io_op_bits_active_vamo ? _T_2314 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2314 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4797) : _T_4797;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4824 = io_op_bits_active_vamo ? _T_2315 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2315 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4799) : _T_4799;	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4825 = io_op_bits_active_vamo ? _T_2299 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2299 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4786) : _T_4786;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4826 = io_op_bits_active_vamo ? _T_2300 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2300 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4788) : _T_4788;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4827 = io_op_bits_active_vamo ? _T_2301 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2301 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4790) : _T_4790;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4828 = io_op_bits_active_vamo ? _T_2302 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2302 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4792) : _T_4792;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4829 = io_op_bits_active_vamo ? _T_2303 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2303 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4794) : _T_4794;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4830 = io_op_bits_active_vamo ? _T_2304 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2304 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4796) : _T_4796;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4831 = io_op_bits_active_vamo ? _T_2305 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2305 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4798) : _T_4798;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4832 = io_op_bits_active_vamo ? _T_2306 & &_T_2 | ~(&_T_2) & ~(&_T_1) & (_T_2306 & &_T_0 |
                ~(&_T_0) & ~(&tail) & _T_4800) : _T_4800;	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4833 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2279 & &tail | _T_2238 & &tail |
                ~(&tail) & _T_4809) : _T_4809;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4834 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2280 & &tail | _T_2242 & &tail |
                ~(&tail) & _T_4810) : _T_4810;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4835 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2281 & &tail | _T_2246 & &tail |
                ~(&tail) & _T_4811) : _T_4811;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4836 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2282 & &tail | _T_2250 & &tail |
                ~(&tail) & _T_4812) : _T_4812;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4837 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2283 & &tail | _T_2254 & &tail |
                ~(&tail) & _T_4813) : _T_4813;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4838 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2284 & &tail | _T_2258 & &tail |
                ~(&tail) & _T_4814) : _T_4814;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4839 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2285 & &tail | _T_2262 & &tail |
                ~(&tail) & _T_4815) : _T_4815;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4840 = io_op_bits_active_vldx ? ~(&_T_1) & ~(&_T_0) & (_T_2286 & &tail | _T_2266 & &tail |
                ~(&tail) & _T_4816) : _T_4816;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4841 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2308 & &_T_1 | ~(&_T_1) & (_T_2308 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4817) : _T_4817);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4842 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2299 & &_T_1 | ~(&_T_1) & (_T_2299 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4825) : _T_4825);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4843 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2309 & &_T_1 | ~(&_T_1) & (_T_2309 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4818) : _T_4818);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4844 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2300 & &_T_1 | ~(&_T_1) & (_T_2300 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4826) : _T_4826);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4845 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2310 & &_T_1 | ~(&_T_1) & (_T_2310 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4819) : _T_4819);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4846 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2301 & &_T_1 | ~(&_T_1) & (_T_2301 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4827) : _T_4827);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4847 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2311 & &_T_1 | ~(&_T_1) & (_T_2311 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4820) : _T_4820);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4848 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2302 & &_T_1 | ~(&_T_1) & (_T_2302 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4828) : _T_4828);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4849 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2312 & &_T_1 | ~(&_T_1) & (_T_2312 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4821) : _T_4821);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4850 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2303 & &_T_1 | ~(&_T_1) & (_T_2303 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4829) : _T_4829);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4851 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2313 & &_T_1 | ~(&_T_1) & (_T_2313 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4822) : _T_4822);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4852 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2304 & &_T_1 | ~(&_T_1) & (_T_2304 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4830) : _T_4830);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4853 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2314 & &_T_1 | ~(&_T_1) & (_T_2314 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4823) : _T_4823);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4854 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2305 & &_T_1 | ~(&_T_1) & (_T_2305 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4831) : _T_4831);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4855 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2315 & &_T_1 | ~(&_T_1) & (_T_2315 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4824) : _T_4824);	// sequencer-master.scala:132:52, :184:52, :267:35, util.scala:94:11
      wire _T_4856 = (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vldx ?
                _T_2306 & &_T_1 | ~(&_T_1) & (_T_2306 & &_T_0 | ~(&_T_0) & ~(&tail) & _T_4832) : _T_4832);	// sequencer-master.scala:133:52, :185:52, :267:35, util.scala:94:11
      wire _T_4857 = io_op_bits_active_vstx ? &_T_1 & _T_132 | _T_2299 & &_T_1 | _T_2238 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2279 & &tail | _T_2238 & &tail | ~(&tail) & _T_4833) : _T_4833;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4858 = io_op_bits_active_vstx ? &_T_1 & _T_133 | _T_2300 & &_T_1 | _T_2242 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2280 & &tail | _T_2242 & &tail | ~(&tail) & _T_4834) : _T_4834;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4859 = io_op_bits_active_vstx ? &_T_1 & _T_134 | _T_2301 & &_T_1 | _T_2246 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2281 & &tail | _T_2246 & &tail | ~(&tail) & _T_4835) : _T_4835;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4860 = io_op_bits_active_vstx ? &_T_1 & _T_135 | _T_2302 & &_T_1 | _T_2250 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2282 & &tail | _T_2250 & &tail | ~(&tail) & _T_4836) : _T_4836;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4861 = io_op_bits_active_vstx ? &_T_1 & _T_136 | _T_2303 & &_T_1 | _T_2254 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2283 & &tail | _T_2254 & &tail | ~(&tail) & _T_4837) : _T_4837;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4862 = io_op_bits_active_vstx ? &_T_1 & _T_137 | _T_2304 & &_T_1 | _T_2258 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2284 & &tail | _T_2258 & &tail | ~(&tail) & _T_4838) : _T_4838;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4863 = io_op_bits_active_vstx ? &_T_1 & _T_138 | _T_2305 & &_T_1 | _T_2262 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2285 & &tail | _T_2262 & &tail | ~(&tail) & _T_4839) : _T_4839;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4864 = io_op_bits_active_vstx ? &_T_1 & &_T_0 | _T_2306 & &_T_1 | _T_2266 & &_T_1 | ~(&_T_1) &
                ~(&_T_0) & (_T_2286 & &tail | _T_2266 & &tail | ~(&tail) & _T_4840) : _T_4840;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4865 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2238 & &tail | ~(&tail) & _T_4857) :
                _T_4857;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4866 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2242 & &tail | ~(&tail) & _T_4858) :
                _T_4858;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4867 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2246 & &tail | ~(&tail) & _T_4859) :
                _T_4859;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4868 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2250 & &tail | ~(&tail) & _T_4860) :
                _T_4860;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4869 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2254 & &tail | ~(&tail) & _T_4861) :
                _T_4861;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4870 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2258 & &tail | ~(&tail) & _T_4862) :
                _T_4862;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4871 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2262 & &tail | ~(&tail) & _T_4863) :
                _T_4863;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
      wire _T_4872 = io_op_bits_active_vld ? ~(&_T_1) & ~(&_T_0) & (_T_2266 & &tail | ~(&tail) & _T_4864) :
                _T_4864;	// sequencer-master.scala:131:52, :183:52, :267:35, util.scala:94:11
  always @(posedge clock) begin	// sequencer-master.scala:107:14
    `ifndef SYNTHESIS	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2325)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2325)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2326)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2326)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2327)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2327)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2328)	// sequencer-master.scala:298:15, :361:15
        $fwrite(32'h80000002, "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n");	// sequencer-master.scala:298:15
      if (`STOP_COND_ & _T_2328)	// sequencer-master.scala:298:15, :361:15
        $fatal;	// sequencer-master.scala:298:15
      if (`PRINTF_COND_ & _T_2329)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2329)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
    `endif
    if (_T_3) begin	// sequencer-master.scala:332:31
      e_0_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_4 | _T_401 ?
                                                io_op_bits_base_vs3_id : e_0_base_vs3_id) : _T_401 ? io_op_bits_base_vs3_id :
                                                e_0_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_0_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_4 | _T_402 ?
                                                io_op_bits_base_vs3_scalar : e_0_base_vs3_scalar) : _T_402 ? io_op_bits_base_vs3_scalar :
                                                e_0_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_0_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_4 | _T_403 ?
                                                io_op_bits_base_vs3_pred : e_0_base_vs3_pred) : _T_403 ? io_op_bits_base_vs3_pred :
                                                e_0_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_0_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_4 | _T_404 ?
                                                io_op_bits_base_vs3_prec : e_0_base_vs3_prec) : _T_404 ? io_op_bits_base_vs3_prec :
                                                e_0_base_vs3_prec;	// sequencer-master.scala:329:29
      e_1_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_5 | _T_405 ?
                                                io_op_bits_base_vs3_id : e_1_base_vs3_id) : _T_405 ? io_op_bits_base_vs3_id :
                                                e_1_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_1_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_5 | _T_406 ?
                                                io_op_bits_base_vs3_scalar : e_1_base_vs3_scalar) : _T_406 ? io_op_bits_base_vs3_scalar :
                                                e_1_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_1_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_5 | _T_407 ?
                                                io_op_bits_base_vs3_pred : e_1_base_vs3_pred) : _T_407 ? io_op_bits_base_vs3_pred :
                                                e_1_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_1_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_5 | _T_408 ?
                                                io_op_bits_base_vs3_prec : e_1_base_vs3_prec) : _T_408 ? io_op_bits_base_vs3_prec :
                                                e_1_base_vs3_prec;	// sequencer-master.scala:329:29
      e_2_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_6 | _T_409 ?
                                                io_op_bits_base_vs3_id : e_2_base_vs3_id) : _T_409 ? io_op_bits_base_vs3_id :
                                                e_2_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_2_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_6 | _T_410 ?
                                                io_op_bits_base_vs3_scalar : e_2_base_vs3_scalar) : _T_410 ? io_op_bits_base_vs3_scalar :
                                                e_2_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_2_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_6 | _T_411 ?
                                                io_op_bits_base_vs3_pred : e_2_base_vs3_pred) : _T_411 ? io_op_bits_base_vs3_pred :
                                                e_2_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_2_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_6 | _T_412 ?
                                                io_op_bits_base_vs3_prec : e_2_base_vs3_prec) : _T_412 ? io_op_bits_base_vs3_prec :
                                                e_2_base_vs3_prec;	// sequencer-master.scala:329:29
      e_3_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_7 | _T_413 ?
                                                io_op_bits_base_vs3_id : e_3_base_vs3_id) : _T_413 ? io_op_bits_base_vs3_id :
                                                e_3_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_3_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_7 | _T_414 ?
                                                io_op_bits_base_vs3_scalar : e_3_base_vs3_scalar) : _T_414 ? io_op_bits_base_vs3_scalar :
                                                e_3_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_3_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_7 | _T_415 ?
                                                io_op_bits_base_vs3_pred : e_3_base_vs3_pred) : _T_415 ? io_op_bits_base_vs3_pred :
                                                e_3_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_3_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_7 | _T_416 ?
                                                io_op_bits_base_vs3_prec : e_3_base_vs3_prec) : _T_416 ? io_op_bits_base_vs3_prec :
                                                e_3_base_vs3_prec;	// sequencer-master.scala:329:29
      e_4_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_8 | _T_417 ?
                                                io_op_bits_base_vs3_id : e_4_base_vs3_id) : _T_417 ? io_op_bits_base_vs3_id :
                                                e_4_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_4_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_8 | _T_418 ?
                                                io_op_bits_base_vs3_scalar : e_4_base_vs3_scalar) : _T_418 ? io_op_bits_base_vs3_scalar :
                                                e_4_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_4_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_8 | _T_419 ?
                                                io_op_bits_base_vs3_pred : e_4_base_vs3_pred) : _T_419 ? io_op_bits_base_vs3_pred :
                                                e_4_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_4_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_8 | _T_420 ?
                                                io_op_bits_base_vs3_prec : e_4_base_vs3_prec) : _T_420 ? io_op_bits_base_vs3_prec :
                                                e_4_base_vs3_prec;	// sequencer-master.scala:329:29
      e_5_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_9 | _T_421 ?
                                                io_op_bits_base_vs3_id : e_5_base_vs3_id) : _T_421 ? io_op_bits_base_vs3_id :
                                                e_5_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_5_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_9 | _T_422 ?
                                                io_op_bits_base_vs3_scalar : e_5_base_vs3_scalar) : _T_422 ? io_op_bits_base_vs3_scalar :
                                                e_5_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_5_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_9 | _T_423 ?
                                                io_op_bits_base_vs3_pred : e_5_base_vs3_pred) : _T_423 ? io_op_bits_base_vs3_pred :
                                                e_5_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_5_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_9 | _T_424 ?
                                                io_op_bits_base_vs3_prec : e_5_base_vs3_prec) : _T_424 ? io_op_bits_base_vs3_prec :
                                                e_5_base_vs3_prec;	// sequencer-master.scala:329:29
      e_6_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_10 | _T_425 ?
                                                io_op_bits_base_vs3_id : e_6_base_vs3_id) : _T_425 ? io_op_bits_base_vs3_id :
                                                e_6_base_vs3_id;	// sequencer-master.scala:141:29, :329:29
      e_6_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_10 | _T_426 ?
                                                io_op_bits_base_vs3_scalar : e_6_base_vs3_scalar) : _T_426 ? io_op_bits_base_vs3_scalar :
                                                e_6_base_vs3_scalar;	// sequencer-master.scala:329:29, types-vxu.scala:119:37
      e_6_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_10 | _T_427 ?
                                                io_op_bits_base_vs3_pred : e_6_base_vs3_pred) : _T_427 ? io_op_bits_base_vs3_pred :
                                                e_6_base_vs3_pred;	// sequencer-master.scala:329:29, types-vxu.scala:119:31
      e_6_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_10 | _T_428 ?
                                                io_op_bits_base_vs3_prec : e_6_base_vs3_prec) : _T_428 ? io_op_bits_base_vs3_prec :
                                                e_6_base_vs3_prec;	// sequencer-master.scala:329:29
      e_7_base_vs3_id <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (&tail | _T_429 ?
                                                io_op_bits_base_vs3_id : e_7_base_vs3_id) : _T_429 ? io_op_bits_base_vs3_id :
                                                e_7_base_vs3_id;	// sequencer-master.scala:141:29, :267:35, :329:29, util.scala:94:11
      e_7_base_vs3_scalar <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (&tail | _T_430 ?
                                                io_op_bits_base_vs3_scalar : e_7_base_vs3_scalar) : _T_430 ? io_op_bits_base_vs3_scalar :
                                                e_7_base_vs3_scalar;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:37, util.scala:94:11
      e_7_base_vs3_pred <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (&tail | _T_431 ?
                                                io_op_bits_base_vs3_pred : e_7_base_vs3_pred) : _T_431 ? io_op_bits_base_vs3_pred :
                                                e_7_base_vs3_pred;	// sequencer-master.scala:267:35, :329:29, types-vxu.scala:119:31, util.scala:94:11
      e_7_base_vs3_prec <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (&tail | _T_432 ?
                                                io_op_bits_base_vs3_prec : e_7_base_vs3_prec) : _T_432 ? io_op_bits_base_vs3_prec :
                                                e_7_base_vs3_prec;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      e_0_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_4 | _T_2330 ?
                                                io_op_bits_sreg_ss3 : e_0_sreg_ss3) : _T_2330 ? io_op_bits_sreg_ss3 : e_0_sreg_ss3;	// sequencer-master.scala:332:31
      e_1_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_5 | _T_2331 ?
                                                io_op_bits_sreg_ss3 : e_1_sreg_ss3) : _T_2331 ? io_op_bits_sreg_ss3 : e_1_sreg_ss3;	// sequencer-master.scala:332:31
      e_2_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_6 | _T_2332 ?
                                                io_op_bits_sreg_ss3 : e_2_sreg_ss3) : _T_2332 ? io_op_bits_sreg_ss3 : e_2_sreg_ss3;	// sequencer-master.scala:332:31
      e_3_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_7 | _T_2333 ?
                                                io_op_bits_sreg_ss3 : e_3_sreg_ss3) : _T_2333 ? io_op_bits_sreg_ss3 : e_3_sreg_ss3;	// sequencer-master.scala:332:31
      e_4_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_8 | _T_2334 ?
                                                io_op_bits_sreg_ss3 : e_4_sreg_ss3) : _T_2334 ? io_op_bits_sreg_ss3 : e_4_sreg_ss3;	// sequencer-master.scala:332:31
      e_5_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_9 | _T_2335 ?
                                                io_op_bits_sreg_ss3 : e_5_sreg_ss3) : _T_2335 ? io_op_bits_sreg_ss3 : e_5_sreg_ss3;	// sequencer-master.scala:332:31
      e_6_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (_T_10 | _T_2336 ?
                                                io_op_bits_sreg_ss3 : e_6_sreg_ss3) : _T_2336 ? io_op_bits_sreg_ss3 : e_6_sreg_ss3;	// sequencer-master.scala:332:31
      e_7_sreg_ss3 <= io_op_bits_active_vfma & io_op_bits_base_vs3_valid & _T_2287 ? (&tail | _T_2337 ?
                                                io_op_bits_sreg_ss3 : e_7_sreg_ss3) : _T_2337 ? io_op_bits_sreg_ss3 : e_7_sreg_ss3;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
    end
    `ifndef SYNTHESIS	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2338)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2338)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2339)	// sequencer-master.scala:298:15, :361:15
        $fwrite(32'h80000002, "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n");	// sequencer-master.scala:298:15
      if (`STOP_COND_ & _T_2339)	// sequencer-master.scala:298:15, :361:15
        $fatal;	// sequencer-master.scala:298:15
      if (`PRINTF_COND_ & _T_2340)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2340)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
    `endif
    if (_T_3) begin	// sequencer-master.scala:332:31
      e_0_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_562 ?
                                                io_op_bits_base_vs2_id : _T_530) : _T_562 ? io_op_bits_base_vs2_id : _T_530;	// sequencer-master.scala:329:29
      e_0_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_563 ?
                                                io_op_bits_base_vs2_scalar : _T_531) : _T_563 ? io_op_bits_base_vs2_scalar : _T_531;	// sequencer-master.scala:329:29
      e_0_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_564 ?
                                                io_op_bits_base_vs2_pred : _T_532) : _T_564 ? io_op_bits_base_vs2_pred : _T_532;	// sequencer-master.scala:329:29
      e_0_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_565 ?
                                                io_op_bits_base_vs2_prec : _T_533) : _T_565 ? io_op_bits_base_vs2_prec : _T_533;	// sequencer-master.scala:329:29
      e_1_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_566 ?
                                                io_op_bits_base_vs2_id : _T_534) : _T_566 ? io_op_bits_base_vs2_id : _T_534;	// sequencer-master.scala:329:29
      e_1_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_567 ?
                                                io_op_bits_base_vs2_scalar : _T_535) : _T_567 ? io_op_bits_base_vs2_scalar : _T_535;	// sequencer-master.scala:329:29
      e_1_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_568 ?
                                                io_op_bits_base_vs2_pred : _T_536) : _T_568 ? io_op_bits_base_vs2_pred : _T_536;	// sequencer-master.scala:329:29
      e_1_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_569 ?
                                                io_op_bits_base_vs2_prec : _T_537) : _T_569 ? io_op_bits_base_vs2_prec : _T_537;	// sequencer-master.scala:329:29
      e_2_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_570 ?
                                                io_op_bits_base_vs2_id : _T_538) : _T_570 ? io_op_bits_base_vs2_id : _T_538;	// sequencer-master.scala:329:29
      e_2_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_571 ?
                                                io_op_bits_base_vs2_scalar : _T_539) : _T_571 ? io_op_bits_base_vs2_scalar : _T_539;	// sequencer-master.scala:329:29
      e_2_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_572 ?
                                                io_op_bits_base_vs2_pred : _T_540) : _T_572 ? io_op_bits_base_vs2_pred : _T_540;	// sequencer-master.scala:329:29
      e_2_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_573 ?
                                                io_op_bits_base_vs2_prec : _T_541) : _T_573 ? io_op_bits_base_vs2_prec : _T_541;	// sequencer-master.scala:329:29
      e_3_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_574 ?
                                                io_op_bits_base_vs2_id : _T_542) : _T_574 ? io_op_bits_base_vs2_id : _T_542;	// sequencer-master.scala:329:29
      e_3_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_575 ?
                                                io_op_bits_base_vs2_scalar : _T_543) : _T_575 ? io_op_bits_base_vs2_scalar : _T_543;	// sequencer-master.scala:329:29
      e_3_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_576 ?
                                                io_op_bits_base_vs2_pred : _T_544) : _T_576 ? io_op_bits_base_vs2_pred : _T_544;	// sequencer-master.scala:329:29
      e_3_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_577 ?
                                                io_op_bits_base_vs2_prec : _T_545) : _T_577 ? io_op_bits_base_vs2_prec : _T_545;	// sequencer-master.scala:329:29
      e_4_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_578 ?
                                                io_op_bits_base_vs2_id : _T_546) : _T_578 ? io_op_bits_base_vs2_id : _T_546;	// sequencer-master.scala:329:29
      e_4_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_579 ?
                                                io_op_bits_base_vs2_scalar : _T_547) : _T_579 ? io_op_bits_base_vs2_scalar : _T_547;	// sequencer-master.scala:329:29
      e_4_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_580 ?
                                                io_op_bits_base_vs2_pred : _T_548) : _T_580 ? io_op_bits_base_vs2_pred : _T_548;	// sequencer-master.scala:329:29
      e_4_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_581 ?
                                                io_op_bits_base_vs2_prec : _T_549) : _T_581 ? io_op_bits_base_vs2_prec : _T_549;	// sequencer-master.scala:329:29
      e_5_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_582 ?
                                                io_op_bits_base_vs2_id : _T_550) : _T_582 ? io_op_bits_base_vs2_id : _T_550;	// sequencer-master.scala:329:29
      e_5_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_583 ?
                                                io_op_bits_base_vs2_scalar : _T_551) : _T_583 ? io_op_bits_base_vs2_scalar : _T_551;	// sequencer-master.scala:329:29
      e_5_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_584 ?
                                                io_op_bits_base_vs2_pred : _T_552) : _T_584 ? io_op_bits_base_vs2_pred : _T_552;	// sequencer-master.scala:329:29
      e_5_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_585 ?
                                                io_op_bits_base_vs2_prec : _T_553) : _T_585 ? io_op_bits_base_vs2_prec : _T_553;	// sequencer-master.scala:329:29
      e_6_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_586 ?
                                                io_op_bits_base_vs2_id : _T_554) : _T_586 ? io_op_bits_base_vs2_id : _T_554;	// sequencer-master.scala:329:29
      e_6_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_587 ?
                                                io_op_bits_base_vs2_scalar : _T_555) : _T_587 ? io_op_bits_base_vs2_scalar : _T_555;	// sequencer-master.scala:329:29
      e_6_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_588 ?
                                                io_op_bits_base_vs2_pred : _T_556) : _T_588 ? io_op_bits_base_vs2_pred : _T_556;	// sequencer-master.scala:329:29
      e_6_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_589 ?
                                                io_op_bits_base_vs2_prec : _T_557) : _T_589 ? io_op_bits_base_vs2_prec : _T_557;	// sequencer-master.scala:329:29
      e_7_base_vs2_id <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_id :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (&tail | _T_590 ?
                                                io_op_bits_base_vs2_id : _T_558) : _T_590 ? io_op_bits_base_vs2_id : _T_558;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      e_7_base_vs2_scalar <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_scalar :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (&tail | _T_591 ?
                                                io_op_bits_base_vs2_scalar : _T_559) : _T_591 ? io_op_bits_base_vs2_scalar : _T_559;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      e_7_base_vs2_pred <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_pred :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (&tail | _T_592 ?
                                                io_op_bits_base_vs2_pred : _T_560) : _T_592 ? io_op_bits_base_vs2_pred : _T_560;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      e_7_base_vs2_prec <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_prec :
                                                io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (&tail | _T_593 ?
                                                io_op_bits_base_vs2_prec : _T_561) : _T_593 ? io_op_bits_base_vs2_prec : _T_561;	// sequencer-master.scala:267:35, :329:29, util.scala:94:11
      e_0_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_4 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_4 | _T_2373 ?
                                                io_op_bits_sreg_ss2 : _T_2365) : _T_2373 ? io_op_bits_sreg_ss2 : _T_2365;	// sequencer-master.scala:332:31
      e_1_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_5 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_5 | _T_2374 ?
                                                io_op_bits_sreg_ss2 : _T_2366) : _T_2374 ? io_op_bits_sreg_ss2 : _T_2366;	// sequencer-master.scala:332:31
      e_2_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_6 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_6 | _T_2375 ?
                                                io_op_bits_sreg_ss2 : _T_2367) : _T_2375 ? io_op_bits_sreg_ss2 : _T_2367;	// sequencer-master.scala:332:31
      e_3_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_7 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_7 | _T_2376 ?
                                                io_op_bits_sreg_ss2 : _T_2368) : _T_2376 ? io_op_bits_sreg_ss2 : _T_2368;	// sequencer-master.scala:332:31
      e_4_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_8 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_8 | _T_2377 ?
                                                io_op_bits_sreg_ss2 : _T_2369) : _T_2377 ? io_op_bits_sreg_ss2 : _T_2369;	// sequencer-master.scala:332:31
      e_5_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_9 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_9 | _T_2378 ?
                                                io_op_bits_sreg_ss2 : _T_2370) : _T_2378 ? io_op_bits_sreg_ss2 : _T_2370;	// sequencer-master.scala:332:31
      e_6_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & _T_10 ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (_T_10 | _T_2379 ?
                                                io_op_bits_sreg_ss2 : _T_2371) : _T_2379 ? io_op_bits_sreg_ss2 : _T_2371;	// sequencer-master.scala:332:31
      e_7_sreg_ss2 <= io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_2277 & &tail ? io_op_bits_sreg_ss2
                                                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid & _T_2277 ? (&tail | _T_2380 ?
                                                io_op_bits_sreg_ss2 : _T_2372) : _T_2380 ? io_op_bits_sreg_ss2 : _T_2372;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
    end
    `ifndef SYNTHESIS	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2381)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2381)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2382)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2382)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2383)	// sequencer-master.scala:298:15, :361:15
        $fwrite(32'h80000002, "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n");	// sequencer-master.scala:298:15
      if (`STOP_COND_ & _T_2383)	// sequencer-master.scala:298:15, :361:15
        $fatal;	// sequencer-master.scala:298:15
      if (`PRINTF_COND_ & _T_2384)	// sequencer-master.scala:298:15, :361:15
        $fwrite(32'h80000002, "Assertion failed: vqu should only be issued for idiv/fdiv/rpred/rfirst\n    at sequencer-master.scala:298 assert(d.active.vidiv || d.active.vfdiv || d.active.vrpred || d.active.vrfirst,\n");	// sequencer-master.scala:298:15
      if (`STOP_COND_ & _T_2384)	// sequencer-master.scala:298:15, :361:15
        $fatal;	// sequencer-master.scala:298:15
      if (`PRINTF_COND_ & _T_2385)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2385)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
      if (`PRINTF_COND_ & _T_2386)	// sequencer-master.scala:361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2386)	// sequencer-master.scala:361:15
        $fatal;	// sequencer-master.scala:361:15
    `endif
    if (_T_3) begin	// sequencer-master.scala:332:31
      e_0_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_4 | _T_2475 ?
                                                io_op_bits_sreg_ss2 : _T_2467) : _T_2475 ? io_op_bits_sreg_ss2 : _T_2467;	// sequencer-master.scala:332:31
      e_1_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_5 | _T_2476 ?
                                                io_op_bits_sreg_ss2 : _T_2468) : _T_2476 ? io_op_bits_sreg_ss2 : _T_2468;	// sequencer-master.scala:332:31
      e_2_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_6 | _T_2477 ?
                                                io_op_bits_sreg_ss2 : _T_2469) : _T_2477 ? io_op_bits_sreg_ss2 : _T_2469;	// sequencer-master.scala:332:31
      e_3_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_7 | _T_2478 ?
                                                io_op_bits_sreg_ss2 : _T_2470) : _T_2478 ? io_op_bits_sreg_ss2 : _T_2470;	// sequencer-master.scala:332:31
      e_4_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_8 | _T_2479 ?
                                                io_op_bits_sreg_ss2 : _T_2471) : _T_2479 ? io_op_bits_sreg_ss2 : _T_2471;	// sequencer-master.scala:332:31
      e_5_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_9 | _T_2480 ?
                                                io_op_bits_sreg_ss2 : _T_2472) : _T_2480 ? io_op_bits_sreg_ss2 : _T_2472;	// sequencer-master.scala:332:31
      e_6_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (_T_10 | _T_2481 ?
                                                io_op_bits_sreg_ss2 : _T_2473) : _T_2481 ? io_op_bits_sreg_ss2 : _T_2473;	// sequencer-master.scala:332:31
      e_7_sreg_ss1 <= io_op_bits_active_vstx & io_op_bits_base_vs2_valid & _T_2277 ? (&tail | _T_2482 ?
                                                io_op_bits_sreg_ss2 : _T_2474) : _T_2482 ? io_op_bits_sreg_ss2 : _T_2474;	// sequencer-master.scala:267:35, :332:31, util.scala:94:11
    end
    `ifndef SYNTHESIS	// sequencer-master.scala:353:15
      if (`PRINTF_COND_ & _T_2483)	// sequencer-master.scala:353:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd_as_vs1: vd should always be vector\n    at sequencer-master.scala:353 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd_as_vs1: vd should always be vector\")\n");	// sequencer-master.scala:353:15
      if (`STOP_COND_ & _T_2483)	// sequencer-master.scala:353:15
        $fatal;	// sequencer-master.scala:353:15
      if (`PRINTF_COND_ & _T_2484)	// sequencer-master.scala:353:15, :361:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd: vd should always be vector\n    at sequencer-master.scala:361 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd: vd should always be vector\")\n");	// sequencer-master.scala:361:15
      if (`STOP_COND_ & _T_2484)	// sequencer-master.scala:353:15, :361:15
        $fatal;	// sequencer-master.scala:361:15
    `endif
    if (_T_3) begin	// sequencer-master.scala:321:24
      e_0_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_291 | _T_1383 ?
                                                io_op_bits_base_vd_id : _T_1205) : _T_1383 ? io_op_bits_base_vd_id : _T_1205;	// sequencer-master.scala:363:24
      e_0_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_291 | _T_1385 ?
                                                io_op_bits_base_vd_scalar : _T_1206) : _T_1385 ? io_op_bits_base_vd_scalar : _T_1206;	// sequencer-master.scala:363:24
      e_0_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_291 | _T_1386 ?
                                                io_op_bits_base_vd_pred : _T_1207) : _T_1386 ? io_op_bits_base_vd_pred : _T_1207;	// sequencer-master.scala:363:24
      e_0_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_291 | _T_1387 ?
                                                io_op_bits_base_vd_prec : _T_1208) : _T_1387 ? io_op_bits_base_vd_prec : _T_1208;	// sequencer-master.scala:363:24
      e_1_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_292 | _T_1388 ?
                                                io_op_bits_base_vd_id : _T_1209) : _T_1388 ? io_op_bits_base_vd_id : _T_1209;	// sequencer-master.scala:363:24
      e_1_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_292 | _T_1390 ?
                                                io_op_bits_base_vd_scalar : _T_1210) : _T_1390 ? io_op_bits_base_vd_scalar : _T_1210;	// sequencer-master.scala:363:24
      e_1_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_292 | _T_1391 ?
                                                io_op_bits_base_vd_pred : _T_1211) : _T_1391 ? io_op_bits_base_vd_pred : _T_1211;	// sequencer-master.scala:363:24
      e_1_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_292 | _T_1392 ?
                                                io_op_bits_base_vd_prec : _T_1212) : _T_1392 ? io_op_bits_base_vd_prec : _T_1212;	// sequencer-master.scala:363:24
      e_2_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_293 | _T_1393 ?
                                                io_op_bits_base_vd_id : _T_1213) : _T_1393 ? io_op_bits_base_vd_id : _T_1213;	// sequencer-master.scala:363:24
      e_2_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_293 | _T_1395 ?
                                                io_op_bits_base_vd_scalar : _T_1214) : _T_1395 ? io_op_bits_base_vd_scalar : _T_1214;	// sequencer-master.scala:363:24
      e_2_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_293 | _T_1396 ?
                                                io_op_bits_base_vd_pred : _T_1215) : _T_1396 ? io_op_bits_base_vd_pred : _T_1215;	// sequencer-master.scala:363:24
      e_2_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_293 | _T_1397 ?
                                                io_op_bits_base_vd_prec : _T_1216) : _T_1397 ? io_op_bits_base_vd_prec : _T_1216;	// sequencer-master.scala:363:24
      e_3_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_294 | _T_1398 ?
                                                io_op_bits_base_vd_id : _T_1217) : _T_1398 ? io_op_bits_base_vd_id : _T_1217;	// sequencer-master.scala:363:24
      e_3_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_294 | _T_1400 ?
                                                io_op_bits_base_vd_scalar : _T_1218) : _T_1400 ? io_op_bits_base_vd_scalar : _T_1218;	// sequencer-master.scala:363:24
      e_3_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_294 | _T_1401 ?
                                                io_op_bits_base_vd_pred : _T_1219) : _T_1401 ? io_op_bits_base_vd_pred : _T_1219;	// sequencer-master.scala:363:24
      e_3_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_294 | _T_1402 ?
                                                io_op_bits_base_vd_prec : _T_1220) : _T_1402 ? io_op_bits_base_vd_prec : _T_1220;	// sequencer-master.scala:363:24
      e_4_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_295 | _T_1403 ?
                                                io_op_bits_base_vd_id : _T_1221) : _T_1403 ? io_op_bits_base_vd_id : _T_1221;	// sequencer-master.scala:363:24
      e_4_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_295 | _T_1405 ?
                                                io_op_bits_base_vd_scalar : _T_1222) : _T_1405 ? io_op_bits_base_vd_scalar : _T_1222;	// sequencer-master.scala:363:24
      e_4_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_295 | _T_1406 ?
                                                io_op_bits_base_vd_pred : _T_1223) : _T_1406 ? io_op_bits_base_vd_pred : _T_1223;	// sequencer-master.scala:363:24
      e_4_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_295 | _T_1407 ?
                                                io_op_bits_base_vd_prec : _T_1224) : _T_1407 ? io_op_bits_base_vd_prec : _T_1224;	// sequencer-master.scala:363:24
      e_5_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_296 | _T_1408 ?
                                                io_op_bits_base_vd_id : _T_1225) : _T_1408 ? io_op_bits_base_vd_id : _T_1225;	// sequencer-master.scala:363:24
      e_5_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_296 | _T_1410 ?
                                                io_op_bits_base_vd_scalar : _T_1226) : _T_1410 ? io_op_bits_base_vd_scalar : _T_1226;	// sequencer-master.scala:363:24
      e_5_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_296 | _T_1411 ?
                                                io_op_bits_base_vd_pred : _T_1227) : _T_1411 ? io_op_bits_base_vd_pred : _T_1227;	// sequencer-master.scala:363:24
      e_5_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_296 | _T_1412 ?
                                                io_op_bits_base_vd_prec : _T_1228) : _T_1412 ? io_op_bits_base_vd_prec : _T_1228;	// sequencer-master.scala:363:24
      e_6_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_297 | _T_1413 ?
                                                io_op_bits_base_vd_id : _T_1229) : _T_1413 ? io_op_bits_base_vd_id : _T_1229;	// sequencer-master.scala:363:24
      e_6_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_297 | _T_1415 ?
                                                io_op_bits_base_vd_scalar : _T_1230) : _T_1415 ? io_op_bits_base_vd_scalar : _T_1230;	// sequencer-master.scala:363:24
      e_6_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_297 | _T_1416 ?
                                                io_op_bits_base_vd_pred : _T_1231) : _T_1416 ? io_op_bits_base_vd_pred : _T_1231;	// sequencer-master.scala:363:24
      e_6_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_297 | _T_1417 ?
                                                io_op_bits_base_vd_prec : _T_1232) : _T_1417 ? io_op_bits_base_vd_prec : _T_1232;	// sequencer-master.scala:363:24
      e_7_base_vd_id <= io_op_bits_active_vld & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (&_T_1 | _T_1418 ?
                                                io_op_bits_base_vd_id : _T_1233) : _T_1418 ? io_op_bits_base_vd_id : _T_1233;	// sequencer-master.scala:267:35, :363:24
      e_7_base_vd_scalar <= io_op_bits_active_vld & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (&_T_1 | _T_1420 ?
                                                io_op_bits_base_vd_scalar : _T_1234) : _T_1420 ? io_op_bits_base_vd_scalar : _T_1234;	// sequencer-master.scala:267:35, :363:24
      e_7_base_vd_pred <= io_op_bits_active_vld & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (&_T_1 | _T_1421 ?
                                                io_op_bits_base_vd_pred : _T_1235) : _T_1421 ? io_op_bits_base_vd_pred : _T_1235;	// sequencer-master.scala:267:35, :363:24
      e_7_base_vd_prec <= io_op_bits_active_vld & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (&_T_1 | _T_1422 ?
                                                io_op_bits_base_vd_prec : _T_1236) : _T_1422 ? io_op_bits_base_vd_prec : _T_1236;	// sequencer-master.scala:267:35, :363:24
      e_0_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vld | ~_T_291 &
                                                ~_T_132 & ~_T_4) & (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (~io_op_bits_active_vldx | ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vamo | ~_T_314
                                                & ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vrfirst | ~_T_4) &
                                                (~io_op_bits_active_vrpred | ~_T_4) & (~io_op_bits_active_vfconv | ~_T_4) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_base_vs2_valid :
                                                ~_T_4 & _T_1037) : _T_1037);	// sequencer-master.scala:274:29, :329:29
      e_1_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vld | ~_T_292 &
                                                ~_T_133 & ~_T_5) & (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (~io_op_bits_active_vldx | ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vamo | ~_T_315
                                                & ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vrfirst | ~_T_5) &
                                                (~io_op_bits_active_vrpred | ~_T_5) & (~io_op_bits_active_vfconv | ~_T_5) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_base_vs2_valid :
                                                ~_T_5 & _T_1038) : _T_1038);	// sequencer-master.scala:274:29, :329:29
      e_2_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vld | ~_T_293 &
                                                ~_T_134 & ~_T_6) & (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (~io_op_bits_active_vldx | ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vamo | ~_T_316
                                                & ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vrfirst | ~_T_6) &
                                                (~io_op_bits_active_vrpred | ~_T_6) & (~io_op_bits_active_vfconv | ~_T_6) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_base_vs2_valid :
                                                ~_T_6 & _T_1039) : _T_1039);	// sequencer-master.scala:274:29, :329:29
      e_3_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vld | ~_T_294 &
                                                ~_T_135 & ~_T_7) & (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (~io_op_bits_active_vldx | ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vamo | ~_T_317
                                                & ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vrfirst | ~_T_7) &
                                                (~io_op_bits_active_vrpred | ~_T_7) & (~io_op_bits_active_vfconv | ~_T_7) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_base_vs2_valid :
                                                ~_T_7 & _T_1040) : _T_1040);	// sequencer-master.scala:274:29, :329:29
      e_4_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vld | ~_T_295 &
                                                ~_T_136 & ~_T_8) & (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (~io_op_bits_active_vldx | ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vamo | ~_T_318
                                                & ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vrfirst | ~_T_8) &
                                                (~io_op_bits_active_vrpred | ~_T_8) & (~io_op_bits_active_vfconv | ~_T_8) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_base_vs2_valid :
                                                ~_T_8 & _T_1041) : _T_1041);	// sequencer-master.scala:274:29, :329:29
      e_5_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vld | ~_T_296 &
                                                ~_T_137 & ~_T_9) & (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (~io_op_bits_active_vldx | ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vamo | ~_T_319
                                                & ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vrfirst | ~_T_9) &
                                                (~io_op_bits_active_vrpred | ~_T_9) & (~io_op_bits_active_vfconv | ~_T_9) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_base_vs2_valid :
                                                ~_T_9 & _T_1042) : _T_1042);	// sequencer-master.scala:274:29, :329:29
      e_6_base_vs2_valid <= (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vld | ~_T_297 &
                                                ~_T_138 & ~_T_10) & (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (~io_op_bits_active_vldx | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vamo | ~_T_320
                                                & ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vrfirst | ~_T_10) &
                                                (~io_op_bits_active_vrpred | ~_T_10) & (~io_op_bits_active_vfconv | ~_T_10) &
                                                (io_op_bits_active_vfcmp ? (io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_base_vs2_valid :
                                                ~_T_10 & _T_1043) : _T_1043);	// sequencer-master.scala:274:29, :329:29
      e_7_base_vs2_valid <= (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vld |
                                                ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) &
                                                ~(&tail)) & (~io_op_bits_active_vldx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (~io_op_bits_active_vamo | ~(&_T_2) & ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                                                (~io_op_bits_active_vfconv | ~(&tail)) & (io_op_bits_active_vfcmp ?
                                                (io_op_bits_base_vs2_valid & &tail ? io_op_bits_base_vs2_valid : ~(&tail) & _T_1044) :
                                                _T_1044);	// sequencer-master.scala:267:35, :274:29, :329:29, util.scala:94:11
      e_0_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vld | ~_T_291 &
                                                ~_T_132 & ~_T_4) & (~io_op_bits_active_vstx | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (~io_op_bits_active_vldx | ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vamo | ~_T_314
                                                & ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vrfirst | ~_T_4) &
                                                (~io_op_bits_active_vrpred | ~_T_4) & (~io_op_bits_active_vfconv | ~_T_4) &
                                                (~io_op_bits_active_vfcmp | ~_T_4) & (~io_op_bits_active_vfdiv | ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_4 ? io_op_bits_base_vs3_valid :
                                                ~_T_4 & _T_868) : _T_868);	// sequencer-master.scala:275:29, :329:29
      e_1_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vld | ~_T_292 &
                                                ~_T_133 & ~_T_5) & (~io_op_bits_active_vstx | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (~io_op_bits_active_vldx | ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vamo | ~_T_315
                                                & ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vrfirst | ~_T_5) &
                                                (~io_op_bits_active_vrpred | ~_T_5) & (~io_op_bits_active_vfconv | ~_T_5) &
                                                (~io_op_bits_active_vfcmp | ~_T_5) & (~io_op_bits_active_vfdiv | ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_5 ? io_op_bits_base_vs3_valid :
                                                ~_T_5 & _T_869) : _T_869);	// sequencer-master.scala:275:29, :329:29
      e_2_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vld | ~_T_293 &
                                                ~_T_134 & ~_T_6) & (~io_op_bits_active_vstx | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (~io_op_bits_active_vldx | ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vamo | ~_T_316
                                                & ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vrfirst | ~_T_6) &
                                                (~io_op_bits_active_vrpred | ~_T_6) & (~io_op_bits_active_vfconv | ~_T_6) &
                                                (~io_op_bits_active_vfcmp | ~_T_6) & (~io_op_bits_active_vfdiv | ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_6 ? io_op_bits_base_vs3_valid :
                                                ~_T_6 & _T_870) : _T_870);	// sequencer-master.scala:275:29, :329:29
      e_3_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vld | ~_T_294 &
                                                ~_T_135 & ~_T_7) & (~io_op_bits_active_vstx | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (~io_op_bits_active_vldx | ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vamo | ~_T_317
                                                & ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vrfirst | ~_T_7) &
                                                (~io_op_bits_active_vrpred | ~_T_7) & (~io_op_bits_active_vfconv | ~_T_7) &
                                                (~io_op_bits_active_vfcmp | ~_T_7) & (~io_op_bits_active_vfdiv | ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_7 ? io_op_bits_base_vs3_valid :
                                                ~_T_7 & _T_871) : _T_871);	// sequencer-master.scala:275:29, :329:29
      e_4_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vld | ~_T_295 &
                                                ~_T_136 & ~_T_8) & (~io_op_bits_active_vstx | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (~io_op_bits_active_vldx | ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vamo | ~_T_318
                                                & ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vrfirst | ~_T_8) &
                                                (~io_op_bits_active_vrpred | ~_T_8) & (~io_op_bits_active_vfconv | ~_T_8) &
                                                (~io_op_bits_active_vfcmp | ~_T_8) & (~io_op_bits_active_vfdiv | ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_8 ? io_op_bits_base_vs3_valid :
                                                ~_T_8 & _T_872) : _T_872);	// sequencer-master.scala:275:29, :329:29
      e_5_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vld | ~_T_296 &
                                                ~_T_137 & ~_T_9) & (~io_op_bits_active_vstx | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (~io_op_bits_active_vldx | ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vamo | ~_T_319
                                                & ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vrfirst | ~_T_9) &
                                                (~io_op_bits_active_vrpred | ~_T_9) & (~io_op_bits_active_vfconv | ~_T_9) &
                                                (~io_op_bits_active_vfcmp | ~_T_9) & (~io_op_bits_active_vfdiv | ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_9 ? io_op_bits_base_vs3_valid :
                                                ~_T_9 & _T_873) : _T_873);	// sequencer-master.scala:275:29, :329:29
      e_6_base_vs3_valid <= (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vld | ~_T_297 &
                                                ~_T_138 & ~_T_10) & (~io_op_bits_active_vstx | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (~io_op_bits_active_vldx | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vamo | ~_T_320
                                                & ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vrfirst | ~_T_10) &
                                                (~io_op_bits_active_vrpred | ~_T_10) & (~io_op_bits_active_vfconv | ~_T_10) &
                                                (~io_op_bits_active_vfcmp | ~_T_10) & (~io_op_bits_active_vfdiv | ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vfma ? (io_op_bits_base_vs3_valid & _T_10 ? io_op_bits_base_vs3_valid :
                                                ~_T_10 & _T_874) : _T_874);	// sequencer-master.scala:275:29, :329:29
      e_7_base_vs3_valid <= (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vld |
                                                ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vstx | ~(&_T_1) & ~(&_T_0) &
                                                ~(&tail)) & (~io_op_bits_active_vldx | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (~io_op_bits_active_vamo | ~(&_T_2) & ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                                                (~io_op_bits_active_vfconv | ~(&tail)) & (~io_op_bits_active_vfcmp | ~(&tail)) &
                                                (~io_op_bits_active_vfdiv | ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vfma ?
                                                (io_op_bits_base_vs3_valid & &tail ? io_op_bits_base_vs3_valid : ~(&tail) & _T_875) :
                                                _T_875);	// sequencer-master.scala:267:35, :275:29, :329:29, util.scala:94:11
      e_0_base_vd_valid <= (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_valid : ~_T_291 & ~_T_132 & ~_T_4 &
                                                _T_1487) : _T_1487);	// sequencer-master.scala:276:28, :363:24
      e_1_base_vd_valid <= (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_valid : ~_T_292 & ~_T_133 & ~_T_5 &
                                                _T_1488) : _T_1488);	// sequencer-master.scala:276:28, :363:24
      e_2_base_vd_valid <= (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_valid : ~_T_293 & ~_T_134 & ~_T_6 &
                                                _T_1489) : _T_1489);	// sequencer-master.scala:276:28, :363:24
      e_3_base_vd_valid <= (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_valid : ~_T_294 & ~_T_135 & ~_T_7 &
                                                _T_1490) : _T_1490);	// sequencer-master.scala:276:28, :363:24
      e_4_base_vd_valid <= (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_valid : ~_T_295 & ~_T_136 & ~_T_8 &
                                                _T_1491) : _T_1491);	// sequencer-master.scala:276:28, :363:24
      e_5_base_vd_valid <= (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_valid : ~_T_296 & ~_T_137 & ~_T_9 &
                                                _T_1492) : _T_1492);	// sequencer-master.scala:276:28, :363:24
      e_6_base_vd_valid <= (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_valid : ~_T_297 & ~_T_138 & ~_T_10
                                                & _T_1493) : _T_1493);	// sequencer-master.scala:276:28, :363:24
      e_7_base_vd_valid <= (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (io_op_bits_active_vld ?
                                                (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_valid : ~(&_T_1) & ~(&_T_0) &
                                                ~(&tail) & _T_1494) : _T_1494);	// sequencer-master.scala:267:35, :276:28, :363:24, util.scala:94:11
      e_0_fn_union <= io_op_bits_active_vst & (_T_291 | _T_132 | _T_4) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_291 | _T_132 | _T_4 | _T_1495 ? io_op_bits_fn_union : _T_1479)
                                                : _T_1495 ? io_op_bits_fn_union : _T_1479;	// sequencer-master.scala:289:23
      e_1_fn_union <= io_op_bits_active_vst & (_T_292 | _T_133 | _T_5) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_292 | _T_133 | _T_5 | _T_1496 ? io_op_bits_fn_union : _T_1480)
                                                : _T_1496 ? io_op_bits_fn_union : _T_1480;	// sequencer-master.scala:289:23
      e_2_fn_union <= io_op_bits_active_vst & (_T_293 | _T_134 | _T_6) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_293 | _T_134 | _T_6 | _T_1497 ? io_op_bits_fn_union : _T_1481)
                                                : _T_1497 ? io_op_bits_fn_union : _T_1481;	// sequencer-master.scala:289:23
      e_3_fn_union <= io_op_bits_active_vst & (_T_294 | _T_135 | _T_7) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_294 | _T_135 | _T_7 | _T_1498 ? io_op_bits_fn_union : _T_1482)
                                                : _T_1498 ? io_op_bits_fn_union : _T_1482;	// sequencer-master.scala:289:23
      e_4_fn_union <= io_op_bits_active_vst & (_T_295 | _T_136 | _T_8) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_295 | _T_136 | _T_8 | _T_1499 ? io_op_bits_fn_union : _T_1483)
                                                : _T_1499 ? io_op_bits_fn_union : _T_1483;	// sequencer-master.scala:289:23
      e_5_fn_union <= io_op_bits_active_vst & (_T_296 | _T_137 | _T_9) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_296 | _T_137 | _T_9 | _T_1500 ? io_op_bits_fn_union : _T_1484)
                                                : _T_1500 ? io_op_bits_fn_union : _T_1484;	// sequencer-master.scala:289:23
      e_6_fn_union <= io_op_bits_active_vst & (_T_297 | _T_138 | _T_10) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (_T_297 | _T_138 | _T_10 | _T_1501 ? io_op_bits_fn_union : _T_1485)
                                                : _T_1501 ? io_op_bits_fn_union : _T_1485;	// sequencer-master.scala:289:23
      e_7_fn_union <= io_op_bits_active_vst & (&_T_1 | &_T_0 | &tail) ? io_op_bits_fn_union :
                                                io_op_bits_active_vld ? (&_T_1 | &_T_0 | &tail | _T_1502 ? io_op_bits_fn_union : _T_1486) :
                                                _T_1502 ? io_op_bits_fn_union : _T_1486;	// sequencer-master.scala:267:35, :289:23, util.scala:94:11
      e_0_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_4 | _T_1535 ? io_op_bits_base_vp_id : _T_1503) : _T_1536) :
                                                _T_1536;	// sequencer-master.scala:321:24
      e_0_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_291 ? io_op_bits_base_vp_valid :
                                                ~_T_291 & ~_T_132 & (io_op_bits_base_vp_valid & _T_4 ? io_op_bits_base_vp_valid : ~_T_4 &
                                                _T_1583)) : _T_1583;	// sequencer-master.scala:272:28, :321:24
      e_0_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_4 | _T_1537 ? io_op_bits_base_vp_scalar : _T_1505) :
                                                _T_1538) : _T_1538;	// sequencer-master.scala:321:24
      e_0_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_4 | _T_1539 ? io_op_bits_base_vp_pred : _T_1506) : _T_1540)
                                                : _T_1540;	// sequencer-master.scala:321:24
      e_1_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_5 | _T_1541 ? io_op_bits_base_vp_id : _T_1507) : _T_1542) :
                                                _T_1542;	// sequencer-master.scala:321:24
      e_1_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_292 ? io_op_bits_base_vp_valid :
                                                ~_T_292 & ~_T_133 & (io_op_bits_base_vp_valid & _T_5 ? io_op_bits_base_vp_valid : ~_T_5 &
                                                _T_1584)) : _T_1584;	// sequencer-master.scala:272:28, :321:24
      e_1_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_5 | _T_1543 ? io_op_bits_base_vp_scalar : _T_1509) :
                                                _T_1544) : _T_1544;	// sequencer-master.scala:321:24
      e_1_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_5 | _T_1545 ? io_op_bits_base_vp_pred : _T_1510) : _T_1546)
                                                : _T_1546;	// sequencer-master.scala:321:24
      e_2_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_6 | _T_1547 ? io_op_bits_base_vp_id : _T_1511) : _T_1548) :
                                                _T_1548;	// sequencer-master.scala:321:24
      e_2_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_293 ? io_op_bits_base_vp_valid :
                                                ~_T_293 & ~_T_134 & (io_op_bits_base_vp_valid & _T_6 ? io_op_bits_base_vp_valid : ~_T_6 &
                                                _T_1585)) : _T_1585;	// sequencer-master.scala:272:28, :321:24
      e_2_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_6 | _T_1549 ? io_op_bits_base_vp_scalar : _T_1513) :
                                                _T_1550) : _T_1550;	// sequencer-master.scala:321:24
      e_2_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_6 | _T_1551 ? io_op_bits_base_vp_pred : _T_1514) : _T_1552)
                                                : _T_1552;	// sequencer-master.scala:321:24
      e_3_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_7 | _T_1553 ? io_op_bits_base_vp_id : _T_1515) : _T_1554) :
                                                _T_1554;	// sequencer-master.scala:321:24
      e_3_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_294 ? io_op_bits_base_vp_valid :
                                                ~_T_294 & ~_T_135 & (io_op_bits_base_vp_valid & _T_7 ? io_op_bits_base_vp_valid : ~_T_7 &
                                                _T_1586)) : _T_1586;	// sequencer-master.scala:272:28, :321:24
      e_3_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_7 | _T_1555 ? io_op_bits_base_vp_scalar : _T_1517) :
                                                _T_1556) : _T_1556;	// sequencer-master.scala:321:24
      e_3_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_7 | _T_1557 ? io_op_bits_base_vp_pred : _T_1518) : _T_1558)
                                                : _T_1558;	// sequencer-master.scala:321:24
      e_4_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_8 | _T_1559 ? io_op_bits_base_vp_id : _T_1519) : _T_1560) :
                                                _T_1560;	// sequencer-master.scala:321:24
      e_4_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_295 ? io_op_bits_base_vp_valid :
                                                ~_T_295 & ~_T_136 & (io_op_bits_base_vp_valid & _T_8 ? io_op_bits_base_vp_valid : ~_T_8 &
                                                _T_1587)) : _T_1587;	// sequencer-master.scala:272:28, :321:24
      e_4_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_8 | _T_1561 ? io_op_bits_base_vp_scalar : _T_1521) :
                                                _T_1562) : _T_1562;	// sequencer-master.scala:321:24
      e_4_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_8 | _T_1563 ? io_op_bits_base_vp_pred : _T_1522) : _T_1564)
                                                : _T_1564;	// sequencer-master.scala:321:24
      e_5_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_9 | _T_1565 ? io_op_bits_base_vp_id : _T_1523) : _T_1566) :
                                                _T_1566;	// sequencer-master.scala:321:24
      e_5_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_296 ? io_op_bits_base_vp_valid :
                                                ~_T_296 & ~_T_137 & (io_op_bits_base_vp_valid & _T_9 ? io_op_bits_base_vp_valid : ~_T_9 &
                                                _T_1588)) : _T_1588;	// sequencer-master.scala:272:28, :321:24
      e_5_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_9 | _T_1567 ? io_op_bits_base_vp_scalar : _T_1525) :
                                                _T_1568) : _T_1568;	// sequencer-master.scala:321:24
      e_5_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_9 | _T_1569 ? io_op_bits_base_vp_pred : _T_1526) : _T_1570)
                                                : _T_1570;	// sequencer-master.scala:321:24
      e_6_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (_T_10 | _T_1571 ? io_op_bits_base_vp_id : _T_1527) : _T_1572) :
                                                _T_1572;	// sequencer-master.scala:321:24
      e_6_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & _T_297 ? io_op_bits_base_vp_valid :
                                                ~_T_297 & ~_T_138 & (io_op_bits_base_vp_valid & _T_10 ? io_op_bits_base_vp_valid : ~_T_10 &
                                                _T_1589)) : _T_1589;	// sequencer-master.scala:272:28, :321:24
      e_6_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (_T_10 | _T_1573 ? io_op_bits_base_vp_scalar : _T_1529) :
                                                _T_1574) : _T_1574;	// sequencer-master.scala:321:24
      e_6_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (_T_10 | _T_1575 ? io_op_bits_base_vp_pred : _T_1530) : _T_1576)
                                                : _T_1576;	// sequencer-master.scala:321:24
      e_7_base_vp_id <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_id :
                                                io_op_bits_base_vp_valid ? (&tail | _T_1577 ? io_op_bits_base_vp_id : _T_1531) : _T_1578) :
                                                _T_1578;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      e_7_base_vp_valid <= io_op_bits_active_vst ? (io_op_bits_base_vp_valid & &_T_1 ? io_op_bits_base_vp_valid :
                                                ~(&_T_1) & ~(&_T_0) & (io_op_bits_base_vp_valid & &tail ? io_op_bits_base_vp_valid :
                                                ~(&tail) & _T_1590)) : _T_1590;	// sequencer-master.scala:267:35, :272:28, :321:24, util.scala:94:11
      e_7_base_vp_scalar <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_scalar :
                                                io_op_bits_base_vp_valid ? (&tail | _T_1579 ? io_op_bits_base_vp_scalar : _T_1533) :
                                                _T_1580) : _T_1580;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
      e_7_base_vp_pred <= io_op_bits_active_vst & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_base_vp_pred :
                                                io_op_bits_base_vp_valid ? (&tail | _T_1581 ? io_op_bits_base_vp_pred : _T_1534) : _T_1582)
                                                : _T_1582;	// sequencer-master.scala:267:35, :321:24, util.scala:94:11
    end
    `ifndef SYNTHESIS	// sequencer-master.scala:353:15
      if (`PRINTF_COND_ & _T_2485)	// sequencer-master.scala:353:15
        $fwrite(32'h80000002, "Assertion failed: iwindow.set.vd_as_vs1: vd should always be vector\n    at sequencer-master.scala:353 assert(!io.op.bits.base.vd.valid || !io.op.bits.base.vd.is_scalar(), \"iwindow.set.vd_as_vs1: vd should always be vector\")\n");	// sequencer-master.scala:353:15
      if (`STOP_COND_ & _T_2485)	// sequencer-master.scala:353:15
        $fatal;	// sequencer-master.scala:353:15
    `endif
    if (_T_3) begin	// sequencer-master.scala:232:25
      e_0_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_4 | _T_2127 ? io_op_bits_base_vs2_id : _T_2071) : _T_2128)
                                                : _T_2128;	// sequencer-master.scala:329:29, :355:25
      e_0_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_valid :
                                                ~_T_291 & ~_T_132 & ~_T_4 & _T_2215) : _T_2215;	// sequencer-master.scala:273:29, :355:25
      e_0_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_4 | _T_2129 ? io_op_bits_base_vs2_scalar : _T_2072) :
                                                _T_2130) : _T_2130;	// sequencer-master.scala:329:29, :355:25
      e_0_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_4 | _T_2131 ? io_op_bits_base_vs2_pred : _T_2073) :
                                                _T_2132) : _T_2132;	// sequencer-master.scala:329:29, :355:25
      e_0_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_4 | _T_2133 ? io_op_bits_base_vs2_prec : _T_2074) :
                                                _T_2134) : _T_2134;	// sequencer-master.scala:329:29, :355:25
      e_1_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_5 | _T_2135 ? io_op_bits_base_vs2_id : _T_2075) : _T_2136)
                                                : _T_2136;	// sequencer-master.scala:329:29, :355:25
      e_1_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_valid :
                                                ~_T_292 & ~_T_133 & ~_T_5 & _T_2216) : _T_2216;	// sequencer-master.scala:273:29, :355:25
      e_1_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_5 | _T_2137 ? io_op_bits_base_vs2_scalar : _T_2076) :
                                                _T_2138) : _T_2138;	// sequencer-master.scala:329:29, :355:25
      e_1_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_5 | _T_2139 ? io_op_bits_base_vs2_pred : _T_2077) :
                                                _T_2140) : _T_2140;	// sequencer-master.scala:329:29, :355:25
      e_1_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_5 | _T_2141 ? io_op_bits_base_vs2_prec : _T_2078) :
                                                _T_2142) : _T_2142;	// sequencer-master.scala:329:29, :355:25
      e_2_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_6 | _T_2143 ? io_op_bits_base_vs2_id : _T_2079) : _T_2144)
                                                : _T_2144;	// sequencer-master.scala:329:29, :355:25
      e_2_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_valid :
                                                ~_T_293 & ~_T_134 & ~_T_6 & _T_2217) : _T_2217;	// sequencer-master.scala:273:29, :355:25
      e_2_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_6 | _T_2145 ? io_op_bits_base_vs2_scalar : _T_2080) :
                                                _T_2146) : _T_2146;	// sequencer-master.scala:329:29, :355:25
      e_2_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_6 | _T_2147 ? io_op_bits_base_vs2_pred : _T_2081) :
                                                _T_2148) : _T_2148;	// sequencer-master.scala:329:29, :355:25
      e_2_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_6 | _T_2149 ? io_op_bits_base_vs2_prec : _T_2082) :
                                                _T_2150) : _T_2150;	// sequencer-master.scala:329:29, :355:25
      e_3_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_7 | _T_2151 ? io_op_bits_base_vs2_id : _T_2083) : _T_2152)
                                                : _T_2152;	// sequencer-master.scala:329:29, :355:25
      e_3_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_valid :
                                                ~_T_294 & ~_T_135 & ~_T_7 & _T_2218) : _T_2218;	// sequencer-master.scala:273:29, :355:25
      e_3_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_7 | _T_2153 ? io_op_bits_base_vs2_scalar : _T_2084) :
                                                _T_2154) : _T_2154;	// sequencer-master.scala:329:29, :355:25
      e_3_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_7 | _T_2155 ? io_op_bits_base_vs2_pred : _T_2085) :
                                                _T_2156) : _T_2156;	// sequencer-master.scala:329:29, :355:25
      e_3_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_7 | _T_2157 ? io_op_bits_base_vs2_prec : _T_2086) :
                                                _T_2158) : _T_2158;	// sequencer-master.scala:329:29, :355:25
      e_4_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_8 | _T_2159 ? io_op_bits_base_vs2_id : _T_2087) : _T_2160)
                                                : _T_2160;	// sequencer-master.scala:329:29, :355:25
      e_4_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_valid :
                                                ~_T_295 & ~_T_136 & ~_T_8 & _T_2219) : _T_2219;	// sequencer-master.scala:273:29, :355:25
      e_4_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_8 | _T_2161 ? io_op_bits_base_vs2_scalar : _T_2088) :
                                                _T_2162) : _T_2162;	// sequencer-master.scala:329:29, :355:25
      e_4_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_8 | _T_2163 ? io_op_bits_base_vs2_pred : _T_2089) :
                                                _T_2164) : _T_2164;	// sequencer-master.scala:329:29, :355:25
      e_4_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_8 | _T_2165 ? io_op_bits_base_vs2_prec : _T_2090) :
                                                _T_2166) : _T_2166;	// sequencer-master.scala:329:29, :355:25
      e_5_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_9 | _T_2167 ? io_op_bits_base_vs2_id : _T_2091) : _T_2168)
                                                : _T_2168;	// sequencer-master.scala:329:29, :355:25
      e_5_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_valid :
                                                ~_T_296 & ~_T_137 & ~_T_9 & _T_2220) : _T_2220;	// sequencer-master.scala:273:29, :355:25
      e_5_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_9 | _T_2169 ? io_op_bits_base_vs2_scalar : _T_2092) :
                                                _T_2170) : _T_2170;	// sequencer-master.scala:329:29, :355:25
      e_5_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_9 | _T_2171 ? io_op_bits_base_vs2_pred : _T_2093) :
                                                _T_2172) : _T_2172;	// sequencer-master.scala:329:29, :355:25
      e_5_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_9 | _T_2173 ? io_op_bits_base_vs2_prec : _T_2094) :
                                                _T_2174) : _T_2174;	// sequencer-master.scala:329:29, :355:25
      e_6_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (_T_10 | _T_2175 ? io_op_bits_base_vs2_id : _T_2095) : _T_2176)
                                                : _T_2176;	// sequencer-master.scala:329:29, :355:25
      e_6_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_valid :
                                                ~_T_297 & ~_T_138 & ~_T_10 & _T_2221) : _T_2221;	// sequencer-master.scala:273:29, :355:25
      e_6_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (_T_10 | _T_2177 ? io_op_bits_base_vs2_scalar : _T_2096) :
                                                _T_2178) : _T_2178;	// sequencer-master.scala:329:29, :355:25
      e_6_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (_T_10 | _T_2179 ? io_op_bits_base_vs2_pred : _T_2097) :
                                                _T_2180) : _T_2180;	// sequencer-master.scala:329:29, :355:25
      e_6_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (_T_10 | _T_2181 ? io_op_bits_base_vs2_prec : _T_2098) :
                                                _T_2182) : _T_2182;	// sequencer-master.scala:329:29, :355:25
      e_7_base_vs1_id <= io_op_bits_active_vst & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_id :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_id :
                                                io_op_bits_base_vs2_valid ? (&tail | _T_2183 ? io_op_bits_base_vs2_id : _T_2099) : _T_2184)
                                                : _T_2184;	// sequencer-master.scala:267:35, :329:29, :355:25, util.scala:94:11
      e_7_base_vs1_valid <= io_op_bits_active_vst ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_valid :
                                                ~(&_T_1) & ~(&_T_0) & ~(&tail) & _T_2222) : _T_2222;	// sequencer-master.scala:267:35, :273:29, :355:25, util.scala:94:11
      e_7_base_vs1_scalar <= io_op_bits_active_vst & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_scalar :
                                                io_op_bits_base_vs2_valid ? (&tail | _T_2185 ? io_op_bits_base_vs2_scalar : _T_2100) :
                                                _T_2186) : _T_2186;	// sequencer-master.scala:267:35, :329:29, :355:25, util.scala:94:11
      e_7_base_vs1_pred <= io_op_bits_active_vst & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_pred :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_pred :
                                                io_op_bits_base_vs2_valid ? (&tail | _T_2187 ? io_op_bits_base_vs2_pred : _T_2101) :
                                                _T_2188) : _T_2188;	// sequencer-master.scala:267:35, :329:29, :355:25, util.scala:94:11
      e_7_base_vs1_prec <= io_op_bits_active_vst & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_prec :
                                                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_base_vd_prec :
                                                io_op_bits_base_vs2_valid ? (&tail | _T_2189 ? io_op_bits_base_vs2_prec : _T_2102) :
                                                _T_2190) : _T_2190;	// sequencer-master.scala:267:35, :329:29, :355:25, util.scala:94:11
      e_0_rports <= io_op_bits_active_vst ? (_T_291 ? _T_2688 : _T_132 | _T_4 | _T_2223 ? 2'h0 : _T_2689) :
                                                _T_2223 ? 2'h0 : _T_2689;	// sequencer-master.scala:230:21, :499:57
      e_1_rports <= io_op_bits_active_vst ? (_T_292 ? _T_2688 : _T_133 | _T_5 | _T_2224 ? 2'h0 : _T_2690) :
                                                _T_2224 ? 2'h0 : _T_2690;	// sequencer-master.scala:230:21, :499:57
      e_2_rports <= io_op_bits_active_vst ? (_T_293 ? _T_2688 : _T_134 | _T_6 | _T_2225 ? 2'h0 : _T_2691) :
                                                _T_2225 ? 2'h0 : _T_2691;	// sequencer-master.scala:230:21, :499:57
      e_3_rports <= io_op_bits_active_vst ? (_T_294 ? _T_2688 : _T_135 | _T_7 | _T_2226 ? 2'h0 : _T_2692) :
                                                _T_2226 ? 2'h0 : _T_2692;	// sequencer-master.scala:230:21, :499:57
      e_4_rports <= io_op_bits_active_vst ? (_T_295 ? _T_2688 : _T_136 | _T_8 | _T_2227 ? 2'h0 : _T_2693) :
                                                _T_2227 ? 2'h0 : _T_2693;	// sequencer-master.scala:230:21, :499:57
      e_5_rports <= io_op_bits_active_vst ? (_T_296 ? _T_2688 : _T_137 | _T_9 | _T_2228 ? 2'h0 : _T_2694) :
                                                _T_2228 ? 2'h0 : _T_2694;	// sequencer-master.scala:230:21, :499:57
      e_6_rports <= io_op_bits_active_vst ? (_T_297 ? _T_2688 : _T_138 | _T_10 | _T_2229 ? 2'h0 : _T_2695) :
                                                _T_2229 ? 2'h0 : _T_2695;	// sequencer-master.scala:230:21, :499:57
      e_7_rports <= io_op_bits_active_vst ? (&_T_1 ? _T_2688 : &_T_0 | &tail | _T_2230 ? 2'h0 : _T_2696) :
                                                _T_2230 ? 2'h0 : _T_2696;	// sequencer-master.scala:230:21, :267:35, :499:57, util.scala:94:11
      e_0_wport_sram <= io_op_bits_active_vst & (_T_291 | _T_132 | _T_4) ? 4'h0 : io_op_bits_active_vld ? (_T_291 |
                                                _T_132 | _T_4 | _T_2199 ? 4'h0 : _T_2672) : _T_2199 ? 4'h0 : _T_2672;	// sequencer-master.scala:231:25, :247:46
      e_1_wport_sram <= io_op_bits_active_vst & (_T_292 | _T_133 | _T_5) ? 4'h0 : io_op_bits_active_vld ? (_T_292 |
                                                _T_133 | _T_5 | _T_2200 ? 4'h0 : _T_2673) : _T_2200 ? 4'h0 : _T_2673;	// sequencer-master.scala:231:25, :247:46
      e_2_wport_sram <= io_op_bits_active_vst & (_T_293 | _T_134 | _T_6) ? 4'h0 : io_op_bits_active_vld ? (_T_293 |
                                                _T_134 | _T_6 | _T_2201 ? 4'h0 : _T_2674) : _T_2201 ? 4'h0 : _T_2674;	// sequencer-master.scala:231:25, :247:46
      e_3_wport_sram <= io_op_bits_active_vst & (_T_294 | _T_135 | _T_7) ? 4'h0 : io_op_bits_active_vld ? (_T_294 |
                                                _T_135 | _T_7 | _T_2202 ? 4'h0 : _T_2675) : _T_2202 ? 4'h0 : _T_2675;	// sequencer-master.scala:231:25, :247:46
      e_4_wport_sram <= io_op_bits_active_vst & (_T_295 | _T_136 | _T_8) ? 4'h0 : io_op_bits_active_vld ? (_T_295 |
                                                _T_136 | _T_8 | _T_2203 ? 4'h0 : _T_2676) : _T_2203 ? 4'h0 : _T_2676;	// sequencer-master.scala:231:25, :247:46
      e_5_wport_sram <= io_op_bits_active_vst & (_T_296 | _T_137 | _T_9) ? 4'h0 : io_op_bits_active_vld ? (_T_296 |
                                                _T_137 | _T_9 | _T_2204 ? 4'h0 : _T_2677) : _T_2204 ? 4'h0 : _T_2677;	// sequencer-master.scala:231:25, :247:46
      e_6_wport_sram <= io_op_bits_active_vst & (_T_297 | _T_138 | _T_10) ? 4'h0 : io_op_bits_active_vld ? (_T_297
                                                | _T_138 | _T_10 | _T_2205 ? 4'h0 : _T_2678) : _T_2205 ? 4'h0 : _T_2678;	// sequencer-master.scala:231:25, :247:46
      e_7_wport_sram <= io_op_bits_active_vst & (&_T_1 | &_T_0 | &tail) ? 4'h0 : io_op_bits_active_vld ? (&_T_1 |
                                                &_T_0 | &tail | _T_2206 ? 4'h0 : _T_2679) : _T_2206 ? 4'h0 : _T_2679;	// sequencer-master.scala:231:25, :247:46, :267:35, util.scala:94:11
      e_0_wport_pred <= io_op_bits_active_vst & (_T_291 | _T_132 | _T_4) ? 3'h0 : io_op_bits_active_vld ? (_T_291 |
                                                _T_132 | _T_4 | _T_2207 ? 3'h0 : _T_2680) : _T_2207 ? 3'h0 : _T_2680;	// sequencer-master.scala:112:17, :232:25
      e_1_wport_pred <= io_op_bits_active_vst & (_T_292 | _T_133 | _T_5) ? 3'h0 : io_op_bits_active_vld ? (_T_292 |
                                                _T_133 | _T_5 | _T_2208 ? 3'h0 : _T_2681) : _T_2208 ? 3'h0 : _T_2681;	// sequencer-master.scala:112:17, :232:25
      e_2_wport_pred <= io_op_bits_active_vst & (_T_293 | _T_134 | _T_6) ? 3'h0 : io_op_bits_active_vld ? (_T_293 |
                                                _T_134 | _T_6 | _T_2209 ? 3'h0 : _T_2682) : _T_2209 ? 3'h0 : _T_2682;	// sequencer-master.scala:112:17, :232:25
      e_3_wport_pred <= io_op_bits_active_vst & (_T_294 | _T_135 | _T_7) ? 3'h0 : io_op_bits_active_vld ? (_T_294 |
                                                _T_135 | _T_7 | _T_2210 ? 3'h0 : _T_2683) : _T_2210 ? 3'h0 : _T_2683;	// sequencer-master.scala:112:17, :232:25
      e_4_wport_pred <= io_op_bits_active_vst & (_T_295 | _T_136 | _T_8) ? 3'h0 : io_op_bits_active_vld ? (_T_295 |
                                                _T_136 | _T_8 | _T_2211 ? 3'h0 : _T_2684) : _T_2211 ? 3'h0 : _T_2684;	// sequencer-master.scala:112:17, :232:25
      e_5_wport_pred <= io_op_bits_active_vst & (_T_296 | _T_137 | _T_9) ? 3'h0 : io_op_bits_active_vld ? (_T_296 |
                                                _T_137 | _T_9 | _T_2212 ? 3'h0 : _T_2685) : _T_2212 ? 3'h0 : _T_2685;	// sequencer-master.scala:112:17, :232:25
      e_6_wport_pred <= io_op_bits_active_vst & (_T_297 | _T_138 | _T_10) ? 3'h0 : io_op_bits_active_vld ? (_T_297
                                                | _T_138 | _T_10 | _T_2213 ? 3'h0 : _T_2686) : _T_2213 ? 3'h0 : _T_2686;	// sequencer-master.scala:112:17, :232:25
      e_7_wport_pred <= io_op_bits_active_vst & (&_T_1 | &_T_0 | &tail) ? 3'h0 : io_op_bits_active_vld ? (&_T_1 |
                                                &_T_0 | &tail | _T_2214 ? 3'h0 : _T_2687) : _T_2214 ? 3'h0 : _T_2687;	// sequencer-master.scala:112:17, :232:25, :267:35, util.scala:94:11
    end
    e_0_last <= io_vf_stop & _T_2317 == 3'h0 | (~_T_3 | (~io_op_bits_active_vst | ~_T_291 & ~_T_132 &
                                ~_T_4) & (~io_op_bits_active_vld | ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vstx |
                                ~_T_291 & ~_T_132 & ~_T_4) & (~io_op_bits_active_vldx | ~_T_291 & ~_T_132 & ~_T_4) &
                                (~io_op_bits_active_vamo | ~_T_314 & ~_T_291 & ~_T_132 & ~_T_4) &
                                (~io_op_bits_active_vrfirst | ~_T_4) & (~io_op_bits_active_vrpred | ~_T_4) &
                                (~io_op_bits_active_vfconv | ~_T_4) & (~io_op_bits_active_vfcmp | ~_T_4) &
                                (~io_op_bits_active_vfdiv | ~_T_132 & ~_T_4) & (~io_op_bits_active_vfma | ~_T_4) &
                                (~io_op_bits_active_vidiv | ~_T_132 & ~_T_4) & (~io_op_bits_active_vimul | ~_T_4) &
                                (~io_op_bits_active_vipred | ~_T_4) & (~io_op_bits_active_vint | ~_T_4)) & e_0_last;	// sequencer-master.scala:112:17, :283:19, :293:19
    e_1_last <= io_vf_stop & _T_2317 == 3'h1 | (~_T_3 | (~io_op_bits_active_vst | ~_T_292 & ~_T_133 &
                                ~_T_5) & (~io_op_bits_active_vld | ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vstx |
                                ~_T_292 & ~_T_133 & ~_T_5) & (~io_op_bits_active_vldx | ~_T_292 & ~_T_133 & ~_T_5) &
                                (~io_op_bits_active_vamo | ~_T_315 & ~_T_292 & ~_T_133 & ~_T_5) &
                                (~io_op_bits_active_vrfirst | ~_T_5) & (~io_op_bits_active_vrpred | ~_T_5) &
                                (~io_op_bits_active_vfconv | ~_T_5) & (~io_op_bits_active_vfcmp | ~_T_5) &
                                (~io_op_bits_active_vfdiv | ~_T_133 & ~_T_5) & (~io_op_bits_active_vfma | ~_T_5) &
                                (~io_op_bits_active_vidiv | ~_T_133 & ~_T_5) & (~io_op_bits_active_vimul | ~_T_5) &
                                (~io_op_bits_active_vipred | ~_T_5) & (~io_op_bits_active_vint | ~_T_5)) & e_1_last;	// sequencer-master.scala:267:35, :283:19, :293:19
    e_2_last <= io_vf_stop & _T_2317 == 3'h2 | (~_T_3 | (~io_op_bits_active_vst | ~_T_293 & ~_T_134 &
                                ~_T_6) & (~io_op_bits_active_vld | ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vstx |
                                ~_T_293 & ~_T_134 & ~_T_6) & (~io_op_bits_active_vldx | ~_T_293 & ~_T_134 & ~_T_6) &
                                (~io_op_bits_active_vamo | ~_T_316 & ~_T_293 & ~_T_134 & ~_T_6) &
                                (~io_op_bits_active_vrfirst | ~_T_6) & (~io_op_bits_active_vrpred | ~_T_6) &
                                (~io_op_bits_active_vfconv | ~_T_6) & (~io_op_bits_active_vfcmp | ~_T_6) &
                                (~io_op_bits_active_vfdiv | ~_T_134 & ~_T_6) & (~io_op_bits_active_vfma | ~_T_6) &
                                (~io_op_bits_active_vidiv | ~_T_134 & ~_T_6) & (~io_op_bits_active_vimul | ~_T_6) &
                                (~io_op_bits_active_vipred | ~_T_6) & (~io_op_bits_active_vint | ~_T_6)) & e_2_last;	// sequencer-master.scala:267:35, :283:19, :293:19
    e_3_last <= io_vf_stop & _T_2317 == 3'h3 | (~_T_3 | (~io_op_bits_active_vst | ~_T_294 & ~_T_135 &
                                ~_T_7) & (~io_op_bits_active_vld | ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vstx |
                                ~_T_294 & ~_T_135 & ~_T_7) & (~io_op_bits_active_vldx | ~_T_294 & ~_T_135 & ~_T_7) &
                                (~io_op_bits_active_vamo | ~_T_317 & ~_T_294 & ~_T_135 & ~_T_7) &
                                (~io_op_bits_active_vrfirst | ~_T_7) & (~io_op_bits_active_vrpred | ~_T_7) &
                                (~io_op_bits_active_vfconv | ~_T_7) & (~io_op_bits_active_vfcmp | ~_T_7) &
                                (~io_op_bits_active_vfdiv | ~_T_135 & ~_T_7) & (~io_op_bits_active_vfma | ~_T_7) &
                                (~io_op_bits_active_vidiv | ~_T_135 & ~_T_7) & (~io_op_bits_active_vimul | ~_T_7) &
                                (~io_op_bits_active_vipred | ~_T_7) & (~io_op_bits_active_vint | ~_T_7)) & e_3_last;	// sequencer-master.scala:267:35, :283:19, :293:19
    e_4_last <= io_vf_stop & _T_2317 == 3'h4 | (~_T_3 | (~io_op_bits_active_vst | ~_T_295 & ~_T_136 &
                                ~_T_8) & (~io_op_bits_active_vld | ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vstx |
                                ~_T_295 & ~_T_136 & ~_T_8) & (~io_op_bits_active_vldx | ~_T_295 & ~_T_136 & ~_T_8) &
                                (~io_op_bits_active_vamo | ~_T_318 & ~_T_295 & ~_T_136 & ~_T_8) &
                                (~io_op_bits_active_vrfirst | ~_T_8) & (~io_op_bits_active_vrpred | ~_T_8) &
                                (~io_op_bits_active_vfconv | ~_T_8) & (~io_op_bits_active_vfcmp | ~_T_8) &
                                (~io_op_bits_active_vfdiv | ~_T_136 & ~_T_8) & (~io_op_bits_active_vfma | ~_T_8) &
                                (~io_op_bits_active_vidiv | ~_T_136 & ~_T_8) & (~io_op_bits_active_vimul | ~_T_8) &
                                (~io_op_bits_active_vipred | ~_T_8) & (~io_op_bits_active_vint | ~_T_8)) & e_4_last;	// sequencer-master.scala:283:19, :293:19, util.scala:94:11
    e_5_last <= io_vf_stop & _T_2317 == 3'h5 | (~_T_3 | (~io_op_bits_active_vst | ~_T_296 & ~_T_137 &
                                ~_T_9) & (~io_op_bits_active_vld | ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vstx |
                                ~_T_296 & ~_T_137 & ~_T_9) & (~io_op_bits_active_vldx | ~_T_296 & ~_T_137 & ~_T_9) &
                                (~io_op_bits_active_vamo | ~_T_319 & ~_T_296 & ~_T_137 & ~_T_9) &
                                (~io_op_bits_active_vrfirst | ~_T_9) & (~io_op_bits_active_vrpred | ~_T_9) &
                                (~io_op_bits_active_vfconv | ~_T_9) & (~io_op_bits_active_vfcmp | ~_T_9) &
                                (~io_op_bits_active_vfdiv | ~_T_137 & ~_T_9) & (~io_op_bits_active_vfma | ~_T_9) &
                                (~io_op_bits_active_vidiv | ~_T_137 & ~_T_9) & (~io_op_bits_active_vimul | ~_T_9) &
                                (~io_op_bits_active_vipred | ~_T_9) & (~io_op_bits_active_vint | ~_T_9)) & e_5_last;	// sequencer-master.scala:183:52, :283:19, :293:19
    e_6_last <= io_vf_stop & _T_2317 == 3'h6 | (~_T_3 | (~io_op_bits_active_vst | ~_T_297 & ~_T_138 &
                                ~_T_10) & (~io_op_bits_active_vld | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vstx
                                | ~_T_297 & ~_T_138 & ~_T_10) & (~io_op_bits_active_vldx | ~_T_297 & ~_T_138 & ~_T_10) &
                                (~io_op_bits_active_vamo | ~_T_320 & ~_T_297 & ~_T_138 & ~_T_10) &
                                (~io_op_bits_active_vrfirst | ~_T_10) & (~io_op_bits_active_vrpred | ~_T_10) &
                                (~io_op_bits_active_vfconv | ~_T_10) & (~io_op_bits_active_vfcmp | ~_T_10) &
                                (~io_op_bits_active_vfdiv | ~_T_138 & ~_T_10) & (~io_op_bits_active_vfma | ~_T_10) &
                                (~io_op_bits_active_vidiv | ~_T_138 & ~_T_10) & (~io_op_bits_active_vimul | ~_T_10) &
                                (~io_op_bits_active_vipred | ~_T_10) & (~io_op_bits_active_vint | ~_T_10)) & e_6_last;	// sequencer-master.scala:267:35, :283:19, :293:19
    e_7_last <= io_vf_stop & &_T_2317 | (~_T_3 | (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail))
                                & (~io_op_bits_active_vld | ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vstx |
                                ~(&_T_1) & ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vldx | ~(&_T_1) & ~(&_T_0) &
                                ~(&tail)) & (~io_op_bits_active_vamo | ~(&_T_2) & ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                (~io_op_bits_active_vrfirst | ~(&tail)) & (~io_op_bits_active_vrpred | ~(&tail)) &
                                (~io_op_bits_active_vfconv | ~(&tail)) & (~io_op_bits_active_vfcmp | ~(&tail)) &
                                (~io_op_bits_active_vfdiv | ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vfma | ~(&tail)) &
                                (~io_op_bits_active_vidiv | ~(&_T_0) & ~(&tail)) & (~io_op_bits_active_vimul | ~(&tail)) &
                                (~io_op_bits_active_vipred | ~(&tail)) & (~io_op_bits_active_vint | ~(&tail))) & e_7_last;	// sequencer-master.scala:267:35, :283:19, :293:19, util.scala:94:11
    _T_2_398 <= _T_397 ? casez_tmp_1 | io_vf_stop & _T_396 == tail : io_vf_stop & ~_T_399;	// sequencer-master.scala:373:43, :435:{17,20}, :441:{17,33,47,58}, :444:24, util.scala:94:11
    if (_T_397 | _T_385) begin	// sequencer-master.scala:188:42, :206:20
      e_0_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_132 | _T_2299 & _T_291
                                                | _T_2238 & _T_291 | ~_T_291 & ~_T_132 & (_T_2238 & _T_4 | ~_T_4 & _T_2961) : _T_2961) :
                                                e_0_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_133 | _T_2300 & _T_291
                                                | _T_2242 & _T_291 | ~_T_291 & ~_T_132 & (_T_2242 & _T_4 | ~_T_4 & _T_2962) : _T_2962) :
                                                e_0_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_134 | _T_2301 & _T_291
                                                | _T_2246 & _T_291 | ~_T_291 & ~_T_132 & (_T_2246 & _T_4 | ~_T_4 & _T_2963) : _T_2963) :
                                                e_0_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_135 | _T_2302 & _T_291
                                                | _T_2250 & _T_291 | ~_T_291 & ~_T_132 & (_T_2250 & _T_4 | ~_T_4 & _T_2964) : _T_2964) :
                                                e_0_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_136 | _T_2303 & _T_291
                                                | _T_2254 & _T_291 | ~_T_291 & ~_T_132 & (_T_2254 & _T_4 | ~_T_4 & _T_2965) : _T_2965) :
                                                e_0_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_137 | _T_2304 & _T_291
                                                | _T_2258 & _T_291 | ~_T_291 & ~_T_132 & (_T_2258 & _T_4 | ~_T_4 & _T_2966) : _T_2966) :
                                                e_0_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & _T_138 | _T_2305 & _T_291
                                                | _T_2262 & _T_291 | ~_T_291 & ~_T_132 & (_T_2262 & _T_4 | ~_T_4 & _T_2967) : _T_2967) :
                                                e_0_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_0_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_291 & &_T_0 | _T_2306 & _T_291 |
                                                _T_2266 & _T_291 | ~_T_291 & ~_T_132 & (_T_2266 & _T_4 | ~_T_4 & _T_2968) : _T_2968) :
                                                e_0_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_0_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_291 | ~_T_291 & (_T_2308 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2937) : _T_2937) : e_0_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_291 | ~_T_291 & (_T_2309 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2939) : _T_2939) : e_0_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_291 | ~_T_291 & (_T_2310 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2941) : _T_2941) : e_0_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_291 | ~_T_291 & (_T_2311 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2943) : _T_2943) : e_0_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_291 | ~_T_291 & (_T_2312 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2945) : _T_2945) : e_0_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_291 | ~_T_291 & (_T_2313 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2947) : _T_2947) : e_0_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_291 | ~_T_291 & (_T_2314 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2949) : _T_2949) : e_0_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_0_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_291 | ~_T_291 & (_T_2315 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2951) : _T_2951) : e_0_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_0_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_291 | ~_T_291 & (_T_2299 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2938) : _T_2938) : e_0_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_291 | ~_T_291 & (_T_2300 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2940) : _T_2940) : e_0_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_291 | ~_T_291 & (_T_2301 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2942) : _T_2942) : e_0_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_291 | ~_T_291 & (_T_2302 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2944) : _T_2944) : e_0_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_291 | ~_T_291 & (_T_2303 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2946) : _T_2946) : e_0_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_291 | ~_T_291 & (_T_2304 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2948) : _T_2948) : e_0_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_291 | ~_T_291 & (_T_2305 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2950) : _T_2950) : e_0_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_0_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_291 & ~_T_132 & ~_T_4) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_291 | ~_T_291 & (_T_2306 & _T_132 | ~_T_132 & ~_T_4 &
                                                _T_2952) : _T_2952) : e_0_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_386) begin	// sequencer-master.scala:188:42, :206:20
      e_1_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_132 | _T_2299 & _T_292
                                                | _T_2238 & _T_292 | ~_T_292 & ~_T_133 & (_T_2238 & _T_5 | ~_T_5 & _T_3233) : _T_3233) :
                                                e_1_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_133 | _T_2300 & _T_292
                                                | _T_2242 & _T_292 | ~_T_292 & ~_T_133 & (_T_2242 & _T_5 | ~_T_5 & _T_3234) : _T_3234) :
                                                e_1_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_134 | _T_2301 & _T_292
                                                | _T_2246 & _T_292 | ~_T_292 & ~_T_133 & (_T_2246 & _T_5 | ~_T_5 & _T_3235) : _T_3235) :
                                                e_1_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_135 | _T_2302 & _T_292
                                                | _T_2250 & _T_292 | ~_T_292 & ~_T_133 & (_T_2250 & _T_5 | ~_T_5 & _T_3236) : _T_3236) :
                                                e_1_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_136 | _T_2303 & _T_292
                                                | _T_2254 & _T_292 | ~_T_292 & ~_T_133 & (_T_2254 & _T_5 | ~_T_5 & _T_3237) : _T_3237) :
                                                e_1_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_137 | _T_2304 & _T_292
                                                | _T_2258 & _T_292 | ~_T_292 & ~_T_133 & (_T_2258 & _T_5 | ~_T_5 & _T_3238) : _T_3238) :
                                                e_1_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & _T_138 | _T_2305 & _T_292
                                                | _T_2262 & _T_292 | ~_T_292 & ~_T_133 & (_T_2262 & _T_5 | ~_T_5 & _T_3239) : _T_3239) :
                                                e_1_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_1_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_292 & &_T_0 | _T_2306 & _T_292 |
                                                _T_2266 & _T_292 | ~_T_292 & ~_T_133 & (_T_2266 & _T_5 | ~_T_5 & _T_3240) : _T_3240) :
                                                e_1_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_1_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_292 | ~_T_292 & (_T_2308 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3209) : _T_3209) : e_1_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_292 | ~_T_292 & (_T_2309 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3211) : _T_3211) : e_1_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_292 | ~_T_292 & (_T_2310 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3213) : _T_3213) : e_1_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_292 | ~_T_292 & (_T_2311 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3215) : _T_3215) : e_1_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_292 | ~_T_292 & (_T_2312 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3217) : _T_3217) : e_1_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_292 | ~_T_292 & (_T_2313 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3219) : _T_3219) : e_1_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_292 | ~_T_292 & (_T_2314 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3221) : _T_3221) : e_1_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_1_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_292 | ~_T_292 & (_T_2315 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3223) : _T_3223) : e_1_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_1_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_292 | ~_T_292 & (_T_2299 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3210) : _T_3210) : e_1_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_292 | ~_T_292 & (_T_2300 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3212) : _T_3212) : e_1_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_292 | ~_T_292 & (_T_2301 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3214) : _T_3214) : e_1_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_292 | ~_T_292 & (_T_2302 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3216) : _T_3216) : e_1_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_292 | ~_T_292 & (_T_2303 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3218) : _T_3218) : e_1_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_292 | ~_T_292 & (_T_2304 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3220) : _T_3220) : e_1_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_292 | ~_T_292 & (_T_2305 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3222) : _T_3222) : e_1_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_1_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_292 & ~_T_133 & ~_T_5) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_292 | ~_T_292 & (_T_2306 & _T_133 | ~_T_133 & ~_T_5 &
                                                _T_3224) : _T_3224) : e_1_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_387) begin	// sequencer-master.scala:188:42, :206:20
      e_2_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_132 | _T_2299 & _T_293
                                                | _T_2238 & _T_293 | ~_T_293 & ~_T_134 & (_T_2238 & _T_6 | ~_T_6 & _T_3505) : _T_3505) :
                                                e_2_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_133 | _T_2300 & _T_293
                                                | _T_2242 & _T_293 | ~_T_293 & ~_T_134 & (_T_2242 & _T_6 | ~_T_6 & _T_3506) : _T_3506) :
                                                e_2_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_134 | _T_2301 & _T_293
                                                | _T_2246 & _T_293 | ~_T_293 & ~_T_134 & (_T_2246 & _T_6 | ~_T_6 & _T_3507) : _T_3507) :
                                                e_2_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_135 | _T_2302 & _T_293
                                                | _T_2250 & _T_293 | ~_T_293 & ~_T_134 & (_T_2250 & _T_6 | ~_T_6 & _T_3508) : _T_3508) :
                                                e_2_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_136 | _T_2303 & _T_293
                                                | _T_2254 & _T_293 | ~_T_293 & ~_T_134 & (_T_2254 & _T_6 | ~_T_6 & _T_3509) : _T_3509) :
                                                e_2_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_137 | _T_2304 & _T_293
                                                | _T_2258 & _T_293 | ~_T_293 & ~_T_134 & (_T_2258 & _T_6 | ~_T_6 & _T_3510) : _T_3510) :
                                                e_2_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & _T_138 | _T_2305 & _T_293
                                                | _T_2262 & _T_293 | ~_T_293 & ~_T_134 & (_T_2262 & _T_6 | ~_T_6 & _T_3511) : _T_3511) :
                                                e_2_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_2_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_293 & &_T_0 | _T_2306 & _T_293 |
                                                _T_2266 & _T_293 | ~_T_293 & ~_T_134 & (_T_2266 & _T_6 | ~_T_6 & _T_3512) : _T_3512) :
                                                e_2_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_2_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_293 | ~_T_293 & (_T_2308 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3481) : _T_3481) : e_2_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_293 | ~_T_293 & (_T_2309 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3483) : _T_3483) : e_2_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_293 | ~_T_293 & (_T_2310 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3485) : _T_3485) : e_2_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_293 | ~_T_293 & (_T_2311 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3487) : _T_3487) : e_2_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_293 | ~_T_293 & (_T_2312 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3489) : _T_3489) : e_2_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_293 | ~_T_293 & (_T_2313 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3491) : _T_3491) : e_2_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_293 | ~_T_293 & (_T_2314 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3493) : _T_3493) : e_2_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_2_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_293 | ~_T_293 & (_T_2315 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3495) : _T_3495) : e_2_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_2_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_293 | ~_T_293 & (_T_2299 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3482) : _T_3482) : e_2_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_293 | ~_T_293 & (_T_2300 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3484) : _T_3484) : e_2_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_293 | ~_T_293 & (_T_2301 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3486) : _T_3486) : e_2_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_293 | ~_T_293 & (_T_2302 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3488) : _T_3488) : e_2_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_293 | ~_T_293 & (_T_2303 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3490) : _T_3490) : e_2_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_293 | ~_T_293 & (_T_2304 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3492) : _T_3492) : e_2_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_293 | ~_T_293 & (_T_2305 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3494) : _T_3494) : e_2_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_2_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_293 & ~_T_134 & ~_T_6) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_293 | ~_T_293 & (_T_2306 & _T_134 | ~_T_134 & ~_T_6 &
                                                _T_3496) : _T_3496) : e_2_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_388) begin	// sequencer-master.scala:188:42, :206:20
      e_3_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_132 | _T_2299 & _T_294
                                                | _T_2238 & _T_294 | ~_T_294 & ~_T_135 & (_T_2238 & _T_7 | ~_T_7 & _T_3777) : _T_3777) :
                                                e_3_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_133 | _T_2300 & _T_294
                                                | _T_2242 & _T_294 | ~_T_294 & ~_T_135 & (_T_2242 & _T_7 | ~_T_7 & _T_3778) : _T_3778) :
                                                e_3_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_134 | _T_2301 & _T_294
                                                | _T_2246 & _T_294 | ~_T_294 & ~_T_135 & (_T_2246 & _T_7 | ~_T_7 & _T_3779) : _T_3779) :
                                                e_3_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_135 | _T_2302 & _T_294
                                                | _T_2250 & _T_294 | ~_T_294 & ~_T_135 & (_T_2250 & _T_7 | ~_T_7 & _T_3780) : _T_3780) :
                                                e_3_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_136 | _T_2303 & _T_294
                                                | _T_2254 & _T_294 | ~_T_294 & ~_T_135 & (_T_2254 & _T_7 | ~_T_7 & _T_3781) : _T_3781) :
                                                e_3_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_137 | _T_2304 & _T_294
                                                | _T_2258 & _T_294 | ~_T_294 & ~_T_135 & (_T_2258 & _T_7 | ~_T_7 & _T_3782) : _T_3782) :
                                                e_3_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & _T_138 | _T_2305 & _T_294
                                                | _T_2262 & _T_294 | ~_T_294 & ~_T_135 & (_T_2262 & _T_7 | ~_T_7 & _T_3783) : _T_3783) :
                                                e_3_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_3_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_294 & &_T_0 | _T_2306 & _T_294 |
                                                _T_2266 & _T_294 | ~_T_294 & ~_T_135 & (_T_2266 & _T_7 | ~_T_7 & _T_3784) : _T_3784) :
                                                e_3_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_3_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_294 | ~_T_294 & (_T_2308 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3753) : _T_3753) : e_3_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_294 | ~_T_294 & (_T_2309 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3755) : _T_3755) : e_3_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_294 | ~_T_294 & (_T_2310 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3757) : _T_3757) : e_3_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_294 | ~_T_294 & (_T_2311 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3759) : _T_3759) : e_3_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_294 | ~_T_294 & (_T_2312 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3761) : _T_3761) : e_3_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_294 | ~_T_294 & (_T_2313 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3763) : _T_3763) : e_3_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_294 | ~_T_294 & (_T_2314 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3765) : _T_3765) : e_3_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_3_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_294 | ~_T_294 & (_T_2315 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3767) : _T_3767) : e_3_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_3_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_294 | ~_T_294 & (_T_2299 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3754) : _T_3754) : e_3_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_294 | ~_T_294 & (_T_2300 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3756) : _T_3756) : e_3_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_294 | ~_T_294 & (_T_2301 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3758) : _T_3758) : e_3_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_294 | ~_T_294 & (_T_2302 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3760) : _T_3760) : e_3_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_294 | ~_T_294 & (_T_2303 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3762) : _T_3762) : e_3_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_294 | ~_T_294 & (_T_2304 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3764) : _T_3764) : e_3_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_294 | ~_T_294 & (_T_2305 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3766) : _T_3766) : e_3_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_3_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_294 & ~_T_135 & ~_T_7) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_294 | ~_T_294 & (_T_2306 & _T_135 | ~_T_135 & ~_T_7 &
                                                _T_3768) : _T_3768) : e_3_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_389) begin	// sequencer-master.scala:188:42, :206:20
      e_4_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_132 | _T_2299 & _T_295
                                                | _T_2238 & _T_295 | ~_T_295 & ~_T_136 & (_T_2238 & _T_8 | ~_T_8 & _T_4049) : _T_4049) :
                                                e_4_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_133 | _T_2300 & _T_295
                                                | _T_2242 & _T_295 | ~_T_295 & ~_T_136 & (_T_2242 & _T_8 | ~_T_8 & _T_4050) : _T_4050) :
                                                e_4_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_134 | _T_2301 & _T_295
                                                | _T_2246 & _T_295 | ~_T_295 & ~_T_136 & (_T_2246 & _T_8 | ~_T_8 & _T_4051) : _T_4051) :
                                                e_4_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_135 | _T_2302 & _T_295
                                                | _T_2250 & _T_295 | ~_T_295 & ~_T_136 & (_T_2250 & _T_8 | ~_T_8 & _T_4052) : _T_4052) :
                                                e_4_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_136 | _T_2303 & _T_295
                                                | _T_2254 & _T_295 | ~_T_295 & ~_T_136 & (_T_2254 & _T_8 | ~_T_8 & _T_4053) : _T_4053) :
                                                e_4_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_137 | _T_2304 & _T_295
                                                | _T_2258 & _T_295 | ~_T_295 & ~_T_136 & (_T_2258 & _T_8 | ~_T_8 & _T_4054) : _T_4054) :
                                                e_4_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & _T_138 | _T_2305 & _T_295
                                                | _T_2262 & _T_295 | ~_T_295 & ~_T_136 & (_T_2262 & _T_8 | ~_T_8 & _T_4055) : _T_4055) :
                                                e_4_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_4_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_295 & &_T_0 | _T_2306 & _T_295 |
                                                _T_2266 & _T_295 | ~_T_295 & ~_T_136 & (_T_2266 & _T_8 | ~_T_8 & _T_4056) : _T_4056) :
                                                e_4_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_4_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_295 | ~_T_295 & (_T_2308 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4025) : _T_4025) : e_4_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_295 | ~_T_295 & (_T_2309 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4027) : _T_4027) : e_4_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_295 | ~_T_295 & (_T_2310 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4029) : _T_4029) : e_4_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_295 | ~_T_295 & (_T_2311 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4031) : _T_4031) : e_4_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_295 | ~_T_295 & (_T_2312 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4033) : _T_4033) : e_4_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_295 | ~_T_295 & (_T_2313 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4035) : _T_4035) : e_4_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_295 | ~_T_295 & (_T_2314 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4037) : _T_4037) : e_4_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_4_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_295 | ~_T_295 & (_T_2315 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4039) : _T_4039) : e_4_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_4_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_295 | ~_T_295 & (_T_2299 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4026) : _T_4026) : e_4_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_295 | ~_T_295 & (_T_2300 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4028) : _T_4028) : e_4_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_295 | ~_T_295 & (_T_2301 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4030) : _T_4030) : e_4_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_295 | ~_T_295 & (_T_2302 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4032) : _T_4032) : e_4_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_295 | ~_T_295 & (_T_2303 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4034) : _T_4034) : e_4_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_295 | ~_T_295 & (_T_2304 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4036) : _T_4036) : e_4_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_295 | ~_T_295 & (_T_2305 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4038) : _T_4038) : e_4_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_4_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_295 & ~_T_136 & ~_T_8) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_295 | ~_T_295 & (_T_2306 & _T_136 | ~_T_136 & ~_T_8 &
                                                _T_4040) : _T_4040) : e_4_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_390) begin	// sequencer-master.scala:188:42, :206:20
      e_5_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_132 | _T_2299 & _T_296
                                                | _T_2238 & _T_296 | ~_T_296 & ~_T_137 & (_T_2238 & _T_9 | ~_T_9 & _T_4321) : _T_4321) :
                                                e_5_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_133 | _T_2300 & _T_296
                                                | _T_2242 & _T_296 | ~_T_296 & ~_T_137 & (_T_2242 & _T_9 | ~_T_9 & _T_4322) : _T_4322) :
                                                e_5_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_134 | _T_2301 & _T_296
                                                | _T_2246 & _T_296 | ~_T_296 & ~_T_137 & (_T_2246 & _T_9 | ~_T_9 & _T_4323) : _T_4323) :
                                                e_5_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_135 | _T_2302 & _T_296
                                                | _T_2250 & _T_296 | ~_T_296 & ~_T_137 & (_T_2250 & _T_9 | ~_T_9 & _T_4324) : _T_4324) :
                                                e_5_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_136 | _T_2303 & _T_296
                                                | _T_2254 & _T_296 | ~_T_296 & ~_T_137 & (_T_2254 & _T_9 | ~_T_9 & _T_4325) : _T_4325) :
                                                e_5_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_137 | _T_2304 & _T_296
                                                | _T_2258 & _T_296 | ~_T_296 & ~_T_137 & (_T_2258 & _T_9 | ~_T_9 & _T_4326) : _T_4326) :
                                                e_5_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & _T_138 | _T_2305 & _T_296
                                                | _T_2262 & _T_296 | ~_T_296 & ~_T_137 & (_T_2262 & _T_9 | ~_T_9 & _T_4327) : _T_4327) :
                                                e_5_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_5_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_296 & &_T_0 | _T_2306 & _T_296 |
                                                _T_2266 & _T_296 | ~_T_296 & ~_T_137 & (_T_2266 & _T_9 | ~_T_9 & _T_4328) : _T_4328) :
                                                e_5_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_5_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_296 | ~_T_296 & (_T_2308 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4297) : _T_4297) : e_5_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_296 | ~_T_296 & (_T_2309 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4299) : _T_4299) : e_5_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_296 | ~_T_296 & (_T_2310 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4301) : _T_4301) : e_5_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_296 | ~_T_296 & (_T_2311 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4303) : _T_4303) : e_5_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_296 | ~_T_296 & (_T_2312 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4305) : _T_4305) : e_5_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_296 | ~_T_296 & (_T_2313 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4307) : _T_4307) : e_5_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_296 | ~_T_296 & (_T_2314 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4309) : _T_4309) : e_5_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_5_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_296 | ~_T_296 & (_T_2315 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4311) : _T_4311) : e_5_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_5_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_296 | ~_T_296 & (_T_2299 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4298) : _T_4298) : e_5_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_296 | ~_T_296 & (_T_2300 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4300) : _T_4300) : e_5_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_296 | ~_T_296 & (_T_2301 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4302) : _T_4302) : e_5_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_296 | ~_T_296 & (_T_2302 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4304) : _T_4304) : e_5_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_296 | ~_T_296 & (_T_2303 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4306) : _T_4306) : e_5_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_296 | ~_T_296 & (_T_2304 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4308) : _T_4308) : e_5_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_296 | ~_T_296 & (_T_2305 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4310) : _T_4310) : e_5_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_5_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_296 & ~_T_137 & ~_T_9) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_296 | ~_T_296 & (_T_2306 & _T_137 | ~_T_137 & ~_T_9 &
                                                _T_4312) : _T_4312) : e_5_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_391) begin	// sequencer-master.scala:188:42, :206:20
      e_6_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_132 | _T_2299 & _T_297
                                                | _T_2238 & _T_297 | ~_T_297 & ~_T_138 & (_T_2238 & _T_10 | ~_T_10 & _T_4593) : _T_4593) :
                                                e_6_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_133 | _T_2300 & _T_297
                                                | _T_2242 & _T_297 | ~_T_297 & ~_T_138 & (_T_2242 & _T_10 | ~_T_10 & _T_4594) : _T_4594) :
                                                e_6_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_134 | _T_2301 & _T_297
                                                | _T_2246 & _T_297 | ~_T_297 & ~_T_138 & (_T_2246 & _T_10 | ~_T_10 & _T_4595) : _T_4595) :
                                                e_6_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_135 | _T_2302 & _T_297
                                                | _T_2250 & _T_297 | ~_T_297 & ~_T_138 & (_T_2250 & _T_10 | ~_T_10 & _T_4596) : _T_4596) :
                                                e_6_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_136 | _T_2303 & _T_297
                                                | _T_2254 & _T_297 | ~_T_297 & ~_T_138 & (_T_2254 & _T_10 | ~_T_10 & _T_4597) : _T_4597) :
                                                e_6_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_137 | _T_2304 & _T_297
                                                | _T_2258 & _T_297 | ~_T_297 & ~_T_138 & (_T_2258 & _T_10 | ~_T_10 & _T_4598) : _T_4598) :
                                                e_6_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & _T_138 | _T_2305 & _T_297
                                                | _T_2262 & _T_297 | ~_T_297 & ~_T_138 & (_T_2262 & _T_10 | ~_T_10 & _T_4599) : _T_4599) :
                                                e_6_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20
      e_6_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? _T_297 & &_T_0 | _T_2306 & _T_297 |
                                                _T_2266 & _T_297 | ~_T_297 & ~_T_138 & (_T_2266 & _T_10 | ~_T_10 & _T_4600) : _T_4600) :
                                                e_6_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21
      e_6_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2308 & _T_297 | ~_T_297 & (_T_2308 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4569) : _T_4569) : e_6_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2309 & _T_297 | ~_T_297 & (_T_2309 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4571) : _T_4571) : e_6_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2310 & _T_297 | ~_T_297 & (_T_2310 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4573) : _T_4573) : e_6_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2311 & _T_297 | ~_T_297 & (_T_2311 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4575) : _T_4575) : e_6_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2312 & _T_297 | ~_T_297 & (_T_2312 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4577) : _T_4577) : e_6_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2313 & _T_297 | ~_T_297 & (_T_2313 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4579) : _T_4579) : e_6_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2314 & _T_297 | ~_T_297 & (_T_2314 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4581) : _T_4581) : e_6_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20
      e_6_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2315 & _T_297 | ~_T_297 & (_T_2315 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4583) : _T_4583) : e_6_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :389:36, :438:21
      e_6_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2299 & _T_297 | ~_T_297 & (_T_2299 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4570) : _T_4570) : e_6_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2300 & _T_297 | ~_T_297 & (_T_2300 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4572) : _T_4572) : e_6_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2301 & _T_297 | ~_T_297 & (_T_2301 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4574) : _T_4574) : e_6_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2302 & _T_297 | ~_T_297 & (_T_2302 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4576) : _T_4576) : e_6_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2303 & _T_297 | ~_T_297 & (_T_2303 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4578) : _T_4578) : e_6_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2304 & _T_297 | ~_T_297 & (_T_2304 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4580) : _T_4580) : e_6_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2305 & _T_297 | ~_T_297 & (_T_2305 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4582) : _T_4582) : e_6_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20
      e_6_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~_T_297 & ~_T_138 & ~_T_10) &
                                                (io_op_bits_active_vld ? _T_2306 & _T_297 | ~_T_297 & (_T_2306 & _T_138 | ~_T_138 & ~_T_10
                                                & _T_4584) : _T_4584) : e_6_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :389:36, :438:21
    end
    if (_T_397 | _T_392) begin	// sequencer-master.scala:188:42, :206:20
      e_7_raw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_132 | _T_2299 & &_T_1 |
                                                _T_2238 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2238 & &tail | ~(&tail) & _T_4865) : _T_4865) :
                                                e_7_raw_0);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_133 | _T_2300 & &_T_1 |
                                                _T_2242 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2242 & &tail | ~(&tail) & _T_4866) : _T_4866) :
                                                e_7_raw_1);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_134 | _T_2301 & &_T_1 |
                                                _T_2246 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2246 & &tail | ~(&tail) & _T_4867) : _T_4867) :
                                                e_7_raw_2);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_135 | _T_2302 & &_T_1 |
                                                _T_2250 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2250 & &tail | ~(&tail) & _T_4868) : _T_4868) :
                                                e_7_raw_3);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_136 | _T_2303 & &_T_1 |
                                                _T_2254 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2254 & &tail | ~(&tail) & _T_4869) : _T_4869) :
                                                e_7_raw_4);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_137 | _T_2304 & &_T_1 |
                                                _T_2258 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2258 & &tail | ~(&tail) & _T_4870) : _T_4870) :
                                                e_7_raw_5);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & _T_138 | _T_2305 & &_T_1 |
                                                _T_2262 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2262 & &tail | ~(&tail) & _T_4871) : _T_4871) :
                                                e_7_raw_6);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, util.scala:94:11
      e_7_raw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (io_op_bits_active_vst ? &_T_1 & &_T_0 | _T_2306 & &_T_1 |
                                                _T_2266 & &_T_1 | ~(&_T_1) & ~(&_T_0) & (_T_2266 & &tail | ~(&tail) & _T_4872) : _T_4872) :
                                                e_7_raw_7);	// sequencer-master.scala:131:52, :183:52, :204:20, :267:35, :389:36, :438:21, util.scala:94:11
      e_7_war_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2308 & &_T_1 | ~(&_T_1) & (_T_2308 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4841) : _T_4841) : e_7_war_0);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2309 & &_T_1 | ~(&_T_1) & (_T_2309 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4843) : _T_4843) : e_7_war_1);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2310 & &_T_1 | ~(&_T_1) & (_T_2310 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4845) : _T_4845) : e_7_war_2);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2311 & &_T_1 | ~(&_T_1) & (_T_2311 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4847) : _T_4847) : e_7_war_3);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2312 & &_T_1 | ~(&_T_1) & (_T_2312 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4849) : _T_4849) : e_7_war_4);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2313 & &_T_1 | ~(&_T_1) & (_T_2313 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4851) : _T_4851) : e_7_war_5);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2314 & &_T_1 | ~(&_T_1) & (_T_2314 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4853) : _T_4853) : e_7_war_6);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, util.scala:94:11
      e_7_war_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2315 & &_T_1 | ~(&_T_1) & (_T_2315 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4855) : _T_4855) : e_7_war_7);	// sequencer-master.scala:132:52, :184:52, :205:20, :267:35, :389:36, :438:21, util.scala:94:11
      e_7_waw_0 <= (~_T_397 | ~_T_2324) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2299 & &_T_1 | ~(&_T_1) & (_T_2299 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4842) : _T_4842) : e_7_waw_0);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_1 <= (~_T_397 | ~_T_2318) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2300 & &_T_1 | ~(&_T_1) & (_T_2300 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4844) : _T_4844) : e_7_waw_1);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_2 <= (~_T_397 | ~_T_2319) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2301 & &_T_1 | ~(&_T_1) & (_T_2301 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4846) : _T_4846) : e_7_waw_2);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_3 <= (~_T_397 | ~_T_2320) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2302 & &_T_1 | ~(&_T_1) & (_T_2302 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4848) : _T_4848) : e_7_waw_3);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_4 <= (~_T_397 | ~_T_2321) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2303 & &_T_1 | ~(&_T_1) & (_T_2303 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4850) : _T_4850) : e_7_waw_4);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_5 <= (~_T_397 | ~_T_2322) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2304 & &_T_1 | ~(&_T_1) & (_T_2304 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4852) : _T_4852) : e_7_waw_5);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_6 <= (~_T_397 | ~_T_2323) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2305 & &_T_1 | ~(&_T_1) & (_T_2305 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4854) : _T_4854) : e_7_waw_6);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, util.scala:94:11
      e_7_waw_7 <= (~_T_397 | ~(&head)) & (_T_3 ? (~io_op_bits_active_vst | ~(&_T_1) & ~(&_T_0) & ~(&tail)) &
                                                (io_op_bits_active_vld ? _T_2306 & &_T_1 | ~(&_T_1) & (_T_2306 & &_T_0 | ~(&_T_0) &
                                                ~(&tail) & _T_4856) : _T_4856) : e_7_waw_7);	// sequencer-master.scala:133:52, :185:52, :206:20, :267:35, :389:36, :438:21, util.scala:94:11
    end
    if (reset) begin	// sequencer-master.scala:107:14
      v_0 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_1 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_2 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_3 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_4 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_5 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_6 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      v_7 <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:107:14
      e_0_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_0_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_1_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_2_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_3_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_4_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_5_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_6_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_viu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vipu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vimu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vidu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vfmu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vfdu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vfcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vfvu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vpu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vgu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vcu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vlu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vsu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      e_7_active_vqu <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:109:14
      maybe_full <= 1'h0;	// compatibility.scala:120:12, sequencer-master.scala:111:23
      head <= 3'h0;	// sequencer-master.scala:112:17
      tail <= 3'h0;	// sequencer-master.scala:112:17, :113:17
    end
    else begin	// sequencer-master.scala:107:14
      tail <= _T_2231 & _T_3 ? (io_op_bits_active_vst | io_op_bits_active_vld | io_op_bits_active_vstx |
                                                io_op_bits_active_vldx ? _T_2 : io_op_bits_active_vamo ? tail - 3'h4 :
                                                io_op_bits_active_vrfirst | io_op_bits_active_vrpred | io_op_bits_active_vfconv |
                                                io_op_bits_active_vfcmp ? _T_0 : io_op_bits_active_vfdiv ? _T_1 : io_op_bits_active_vfma ?
                                                _T_0 : io_op_bits_active_vidiv ? _T_1 : io_op_bits_active_vimul | io_op_bits_active_vipred
                                                | io_op_bits_active_vint ? _T_0 : tail) : tail;	// sequencer-master.scala:265:66, :419:14, util.scala:94:11
      head <= _T_397 ? _T_396 : head;	// sequencer-master.scala:389:36, :423:14
      maybe_full <= ~_T_397 & (_T_2231 | maybe_full);	// sequencer-master.scala:389:15, :420:20, :424:20
      v_0 <= ~reset & (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vst & (_T_291 | _T_132 | _T_4) |
                                                io_op_bits_active_vld & (_T_291 | _T_132 | _T_4) | io_op_bits_active_vstx & (_T_291 |
                                                _T_132 | _T_4) | io_op_bits_active_vldx & (_T_291 | _T_132 | _T_4) | io_op_bits_active_vamo
                                                & (_T_314 | _T_291 | _T_132 | _T_4) | io_op_bits_active_vrfirst & _T_4 |
                                                io_op_bits_active_vrpred & _T_4 | io_op_bits_active_vfconv & _T_4 | io_op_bits_active_vfcmp
                                                & _T_4 | io_op_bits_active_vfdiv & (_T_132 | _T_4) | io_op_bits_active_vfma & _T_4 |
                                                io_op_bits_active_vidiv & (_T_132 | _T_4) | io_op_bits_active_vimul & _T_4 |
                                                io_op_bits_active_vipred & _T_4 | io_op_bits_active_vint & _T_4) | v_0);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_0_active_viu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vint & _T_4 | e_0_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vipu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vipred & _T_4 | e_0_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vimu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vimul & _T_4 | e_0_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vidu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vidiv & _T_132 | e_0_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vfmu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vfma & _T_4 | e_0_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vfdu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vfdiv & _T_132 | e_0_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vfcu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vfcmp & _T_4 | e_0_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vfvu <= (~_T_397 | ~_T_2324) & (_T_3 & io_op_bits_active_vfconv & _T_4 | e_0_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vpu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vst & _T_4 | io_op_bits_active_vld &
                                                _T_4) | e_0_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vgu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vstx & _T_4 | io_op_bits_active_vldx &
                                                _T_4 | io_op_bits_active_vamo & _T_4) | e_0_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vcu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vst & _T_132 | io_op_bits_active_vld &
                                                _T_132 | io_op_bits_active_vstx & _T_132 | io_op_bits_active_vldx & _T_132 |
                                                io_op_bits_active_vamo & _T_132) | e_0_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vlu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vld & _T_291 | io_op_bits_active_vldx &
                                                _T_291 | io_op_bits_active_vamo & _T_314) | e_0_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vsu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vst & _T_291 | io_op_bits_active_vstx &
                                                _T_291 | io_op_bits_active_vamo & _T_291) | e_0_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_0_active_vqu <= (~_T_397 | ~_T_2324) & (_T_3 & (io_op_bits_active_vrfirst & _T_4 | io_op_bits_active_vrpred
                                                & _T_4 | io_op_bits_active_vfdiv & _T_4 | io_op_bits_active_vidiv & _T_4) | e_0_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_1 <= ~reset & (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vst & (_T_292 | _T_133 | _T_5) |
                                                io_op_bits_active_vld & (_T_292 | _T_133 | _T_5) | io_op_bits_active_vstx & (_T_292 |
                                                _T_133 | _T_5) | io_op_bits_active_vldx & (_T_292 | _T_133 | _T_5) | io_op_bits_active_vamo
                                                & (_T_315 | _T_292 | _T_133 | _T_5) | io_op_bits_active_vrfirst & _T_5 |
                                                io_op_bits_active_vrpred & _T_5 | io_op_bits_active_vfconv & _T_5 | io_op_bits_active_vfcmp
                                                & _T_5 | io_op_bits_active_vfdiv & (_T_133 | _T_5) | io_op_bits_active_vfma & _T_5 |
                                                io_op_bits_active_vidiv & (_T_133 | _T_5) | io_op_bits_active_vimul & _T_5 |
                                                io_op_bits_active_vipred & _T_5 | io_op_bits_active_vint & _T_5) | v_1);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_1_active_viu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vint & _T_5 | e_1_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vipu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vipred & _T_5 | e_1_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vimu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vimul & _T_5 | e_1_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vidu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vidiv & _T_133 | e_1_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vfmu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vfma & _T_5 | e_1_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vfdu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vfdiv & _T_133 | e_1_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vfcu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vfcmp & _T_5 | e_1_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vfvu <= (~_T_397 | ~_T_2318) & (_T_3 & io_op_bits_active_vfconv & _T_5 | e_1_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vpu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vst & _T_5 | io_op_bits_active_vld &
                                                _T_5) | e_1_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vgu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vstx & _T_5 | io_op_bits_active_vldx &
                                                _T_5 | io_op_bits_active_vamo & _T_5) | e_1_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vcu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vst & _T_133 | io_op_bits_active_vld &
                                                _T_133 | io_op_bits_active_vstx & _T_133 | io_op_bits_active_vldx & _T_133 |
                                                io_op_bits_active_vamo & _T_133) | e_1_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vlu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vld & _T_292 | io_op_bits_active_vldx &
                                                _T_292 | io_op_bits_active_vamo & _T_315) | e_1_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vsu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vst & _T_292 | io_op_bits_active_vstx &
                                                _T_292 | io_op_bits_active_vamo & _T_292) | e_1_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_1_active_vqu <= (~_T_397 | ~_T_2318) & (_T_3 & (io_op_bits_active_vrfirst & _T_5 | io_op_bits_active_vrpred
                                                & _T_5 | io_op_bits_active_vfdiv & _T_5 | io_op_bits_active_vidiv & _T_5) | e_1_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_2 <= ~reset & (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vst & (_T_293 | _T_134 | _T_6) |
                                                io_op_bits_active_vld & (_T_293 | _T_134 | _T_6) | io_op_bits_active_vstx & (_T_293 |
                                                _T_134 | _T_6) | io_op_bits_active_vldx & (_T_293 | _T_134 | _T_6) | io_op_bits_active_vamo
                                                & (_T_316 | _T_293 | _T_134 | _T_6) | io_op_bits_active_vrfirst & _T_6 |
                                                io_op_bits_active_vrpred & _T_6 | io_op_bits_active_vfconv & _T_6 | io_op_bits_active_vfcmp
                                                & _T_6 | io_op_bits_active_vfdiv & (_T_134 | _T_6) | io_op_bits_active_vfma & _T_6 |
                                                io_op_bits_active_vidiv & (_T_134 | _T_6) | io_op_bits_active_vimul & _T_6 |
                                                io_op_bits_active_vipred & _T_6 | io_op_bits_active_vint & _T_6) | v_2);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_2_active_viu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vint & _T_6 | e_2_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vipu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vipred & _T_6 | e_2_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vimu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vimul & _T_6 | e_2_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vidu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vidiv & _T_134 | e_2_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vfmu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vfma & _T_6 | e_2_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vfdu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vfdiv & _T_134 | e_2_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vfcu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vfcmp & _T_6 | e_2_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vfvu <= (~_T_397 | ~_T_2319) & (_T_3 & io_op_bits_active_vfconv & _T_6 | e_2_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vpu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vst & _T_6 | io_op_bits_active_vld &
                                                _T_6) | e_2_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vgu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vstx & _T_6 | io_op_bits_active_vldx &
                                                _T_6 | io_op_bits_active_vamo & _T_6) | e_2_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vcu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vst & _T_134 | io_op_bits_active_vld &
                                                _T_134 | io_op_bits_active_vstx & _T_134 | io_op_bits_active_vldx & _T_134 |
                                                io_op_bits_active_vamo & _T_134) | e_2_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vlu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vld & _T_293 | io_op_bits_active_vldx &
                                                _T_293 | io_op_bits_active_vamo & _T_316) | e_2_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vsu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vst & _T_293 | io_op_bits_active_vstx &
                                                _T_293 | io_op_bits_active_vamo & _T_293) | e_2_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_2_active_vqu <= (~_T_397 | ~_T_2319) & (_T_3 & (io_op_bits_active_vrfirst & _T_6 | io_op_bits_active_vrpred
                                                & _T_6 | io_op_bits_active_vfdiv & _T_6 | io_op_bits_active_vidiv & _T_6) | e_2_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_3 <= ~reset & (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vst & (_T_294 | _T_135 | _T_7) |
                                                io_op_bits_active_vld & (_T_294 | _T_135 | _T_7) | io_op_bits_active_vstx & (_T_294 |
                                                _T_135 | _T_7) | io_op_bits_active_vldx & (_T_294 | _T_135 | _T_7) | io_op_bits_active_vamo
                                                & (_T_317 | _T_294 | _T_135 | _T_7) | io_op_bits_active_vrfirst & _T_7 |
                                                io_op_bits_active_vrpred & _T_7 | io_op_bits_active_vfconv & _T_7 | io_op_bits_active_vfcmp
                                                & _T_7 | io_op_bits_active_vfdiv & (_T_135 | _T_7) | io_op_bits_active_vfma & _T_7 |
                                                io_op_bits_active_vidiv & (_T_135 | _T_7) | io_op_bits_active_vimul & _T_7 |
                                                io_op_bits_active_vipred & _T_7 | io_op_bits_active_vint & _T_7) | v_3);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_3_active_viu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vint & _T_7 | e_3_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vipu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vipred & _T_7 | e_3_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vimu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vimul & _T_7 | e_3_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vidu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vidiv & _T_135 | e_3_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vfmu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vfma & _T_7 | e_3_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vfdu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vfdiv & _T_135 | e_3_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vfcu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vfcmp & _T_7 | e_3_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vfvu <= (~_T_397 | ~_T_2320) & (_T_3 & io_op_bits_active_vfconv & _T_7 | e_3_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vpu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vst & _T_7 | io_op_bits_active_vld &
                                                _T_7) | e_3_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vgu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vstx & _T_7 | io_op_bits_active_vldx &
                                                _T_7 | io_op_bits_active_vamo & _T_7) | e_3_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vcu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vst & _T_135 | io_op_bits_active_vld &
                                                _T_135 | io_op_bits_active_vstx & _T_135 | io_op_bits_active_vldx & _T_135 |
                                                io_op_bits_active_vamo & _T_135) | e_3_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vlu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vld & _T_294 | io_op_bits_active_vldx &
                                                _T_294 | io_op_bits_active_vamo & _T_317) | e_3_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vsu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vst & _T_294 | io_op_bits_active_vstx &
                                                _T_294 | io_op_bits_active_vamo & _T_294) | e_3_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_3_active_vqu <= (~_T_397 | ~_T_2320) & (_T_3 & (io_op_bits_active_vrfirst & _T_7 | io_op_bits_active_vrpred
                                                & _T_7 | io_op_bits_active_vfdiv & _T_7 | io_op_bits_active_vidiv & _T_7) | e_3_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_4 <= ~reset & (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vst & (_T_295 | _T_136 | _T_8) |
                                                io_op_bits_active_vld & (_T_295 | _T_136 | _T_8) | io_op_bits_active_vstx & (_T_295 |
                                                _T_136 | _T_8) | io_op_bits_active_vldx & (_T_295 | _T_136 | _T_8) | io_op_bits_active_vamo
                                                & (_T_318 | _T_295 | _T_136 | _T_8) | io_op_bits_active_vrfirst & _T_8 |
                                                io_op_bits_active_vrpred & _T_8 | io_op_bits_active_vfconv & _T_8 | io_op_bits_active_vfcmp
                                                & _T_8 | io_op_bits_active_vfdiv & (_T_136 | _T_8) | io_op_bits_active_vfma & _T_8 |
                                                io_op_bits_active_vidiv & (_T_136 | _T_8) | io_op_bits_active_vimul & _T_8 |
                                                io_op_bits_active_vipred & _T_8 | io_op_bits_active_vint & _T_8) | v_4);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_4_active_viu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vint & _T_8 | e_4_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vipu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vipred & _T_8 | e_4_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vimu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vimul & _T_8 | e_4_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vidu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vidiv & _T_136 | e_4_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vfmu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vfma & _T_8 | e_4_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vfdu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vfdiv & _T_136 | e_4_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vfcu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vfcmp & _T_8 | e_4_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vfvu <= (~_T_397 | ~_T_2321) & (_T_3 & io_op_bits_active_vfconv & _T_8 | e_4_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vpu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vst & _T_8 | io_op_bits_active_vld &
                                                _T_8) | e_4_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vgu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vstx & _T_8 | io_op_bits_active_vldx &
                                                _T_8 | io_op_bits_active_vamo & _T_8) | e_4_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vcu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vst & _T_136 | io_op_bits_active_vld &
                                                _T_136 | io_op_bits_active_vstx & _T_136 | io_op_bits_active_vldx & _T_136 |
                                                io_op_bits_active_vamo & _T_136) | e_4_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vlu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vld & _T_295 | io_op_bits_active_vldx &
                                                _T_295 | io_op_bits_active_vamo & _T_318) | e_4_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vsu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vst & _T_295 | io_op_bits_active_vstx &
                                                _T_295 | io_op_bits_active_vamo & _T_295) | e_4_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_4_active_vqu <= (~_T_397 | ~_T_2321) & (_T_3 & (io_op_bits_active_vrfirst & _T_8 | io_op_bits_active_vrpred
                                                & _T_8 | io_op_bits_active_vfdiv & _T_8 | io_op_bits_active_vidiv & _T_8) | e_4_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_5 <= ~reset & (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vst & (_T_296 | _T_137 | _T_9) |
                                                io_op_bits_active_vld & (_T_296 | _T_137 | _T_9) | io_op_bits_active_vstx & (_T_296 |
                                                _T_137 | _T_9) | io_op_bits_active_vldx & (_T_296 | _T_137 | _T_9) | io_op_bits_active_vamo
                                                & (_T_319 | _T_296 | _T_137 | _T_9) | io_op_bits_active_vrfirst & _T_9 |
                                                io_op_bits_active_vrpred & _T_9 | io_op_bits_active_vfconv & _T_9 | io_op_bits_active_vfcmp
                                                & _T_9 | io_op_bits_active_vfdiv & (_T_137 | _T_9) | io_op_bits_active_vfma & _T_9 |
                                                io_op_bits_active_vidiv & (_T_137 | _T_9) | io_op_bits_active_vimul & _T_9 |
                                                io_op_bits_active_vipred & _T_9 | io_op_bits_active_vint & _T_9) | v_5);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_5_active_viu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vint & _T_9 | e_5_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vipu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vipred & _T_9 | e_5_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vimu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vimul & _T_9 | e_5_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vidu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vidiv & _T_137 | e_5_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vfmu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vfma & _T_9 | e_5_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vfdu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vfdiv & _T_137 | e_5_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vfcu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vfcmp & _T_9 | e_5_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vfvu <= (~_T_397 | ~_T_2322) & (_T_3 & io_op_bits_active_vfconv & _T_9 | e_5_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vpu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vst & _T_9 | io_op_bits_active_vld &
                                                _T_9) | e_5_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vgu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vstx & _T_9 | io_op_bits_active_vldx &
                                                _T_9 | io_op_bits_active_vamo & _T_9) | e_5_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vcu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vst & _T_137 | io_op_bits_active_vld &
                                                _T_137 | io_op_bits_active_vstx & _T_137 | io_op_bits_active_vldx & _T_137 |
                                                io_op_bits_active_vamo & _T_137) | e_5_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vlu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vld & _T_296 | io_op_bits_active_vldx &
                                                _T_296 | io_op_bits_active_vamo & _T_319) | e_5_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vsu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vst & _T_296 | io_op_bits_active_vstx &
                                                _T_296 | io_op_bits_active_vamo & _T_296) | e_5_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_5_active_vqu <= (~_T_397 | ~_T_2322) & (_T_3 & (io_op_bits_active_vrfirst & _T_9 | io_op_bits_active_vrpred
                                                & _T_9 | io_op_bits_active_vfdiv & _T_9 | io_op_bits_active_vidiv & _T_9) | e_5_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_6 <= ~reset & (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vst & (_T_297 | _T_138 | _T_10)
                                                | io_op_bits_active_vld & (_T_297 | _T_138 | _T_10) | io_op_bits_active_vstx & (_T_297 |
                                                _T_138 | _T_10) | io_op_bits_active_vldx & (_T_297 | _T_138 | _T_10) |
                                                io_op_bits_active_vamo & (_T_320 | _T_297 | _T_138 | _T_10) | io_op_bits_active_vrfirst &
                                                _T_10 | io_op_bits_active_vrpred & _T_10 | io_op_bits_active_vfconv & _T_10 |
                                                io_op_bits_active_vfcmp & _T_10 | io_op_bits_active_vfdiv & (_T_138 | _T_10) |
                                                io_op_bits_active_vfma & _T_10 | io_op_bits_active_vidiv & (_T_138 | _T_10) |
                                                io_op_bits_active_vimul & _T_10 | io_op_bits_active_vipred & _T_10 | io_op_bits_active_vint
                                                & _T_10) | v_6);	// sequencer-master.scala:136:44, :267:35, :372:35
      e_6_active_viu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vint & _T_10 | e_6_active_viu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vipu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vipred & _T_10 | e_6_active_vipu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vimu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vimul & _T_10 | e_6_active_vimu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vidu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vidiv & _T_138 | e_6_active_vidu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vfmu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vfma & _T_10 | e_6_active_vfmu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vfdu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vfdiv & _T_138 | e_6_active_vfdu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vfcu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vfcmp & _T_10 | e_6_active_vfcu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vfvu <= (~_T_397 | ~_T_2323) & (_T_3 & io_op_bits_active_vfconv & _T_10 | e_6_active_vfvu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vpu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vst & _T_10 | io_op_bits_active_vld &
                                                _T_10) | e_6_active_vpu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vgu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vstx & _T_10 | io_op_bits_active_vldx &
                                                _T_10 | io_op_bits_active_vamo & _T_10) | e_6_active_vgu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vcu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vst & _T_138 | io_op_bits_active_vld &
                                                _T_138 | io_op_bits_active_vstx & _T_138 | io_op_bits_active_vldx & _T_138 |
                                                io_op_bits_active_vamo & _T_138) | e_6_active_vcu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vlu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vld & _T_297 | io_op_bits_active_vldx &
                                                _T_297 | io_op_bits_active_vamo & _T_320) | e_6_active_vlu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vsu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vst & _T_297 | io_op_bits_active_vstx &
                                                _T_297 | io_op_bits_active_vamo & _T_297) | e_6_active_vsu);	// sequencer-master.scala:288:26, :373:43
      e_6_active_vqu <= (~_T_397 | ~_T_2323) & (_T_3 & (io_op_bits_active_vrfirst & _T_10 |
                                                io_op_bits_active_vrpred & _T_10 | io_op_bits_active_vfdiv & _T_10 |
                                                io_op_bits_active_vidiv & _T_10) | e_6_active_vqu);	// sequencer-master.scala:288:26, :373:43
      v_7 <= ~reset & (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vst & (&_T_1 | &_T_0 | &tail) |
                                                io_op_bits_active_vld & (&_T_1 | &_T_0 | &tail) | io_op_bits_active_vstx & (&_T_1 | &_T_0 |
                                                &tail) | io_op_bits_active_vldx & (&_T_1 | &_T_0 | &tail) | io_op_bits_active_vamo & (&_T_2
                                                | &_T_1 | &_T_0 | &tail) | io_op_bits_active_vrfirst & &tail | io_op_bits_active_vrpred &
                                                &tail | io_op_bits_active_vfconv & &tail | io_op_bits_active_vfcmp & &tail |
                                                io_op_bits_active_vfdiv & (&_T_0 | &tail) | io_op_bits_active_vfma & &tail |
                                                io_op_bits_active_vidiv & (&_T_0 | &tail) | io_op_bits_active_vimul & &tail |
                                                io_op_bits_active_vipred & &tail | io_op_bits_active_vint & &tail) | v_7);	// sequencer-master.scala:136:44, :267:35, :372:35, :389:36, :438:21, util.scala:94:11
      e_7_active_viu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vint & &tail | e_7_active_viu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vipu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vipred & &tail | e_7_active_vipu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vimu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vimul & &tail | e_7_active_vimu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vidu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vidiv & &_T_0 | e_7_active_vidu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21
      e_7_active_vfmu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vfma & &tail | e_7_active_vfmu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vfdu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vfdiv & &_T_0 | e_7_active_vfdu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21
      e_7_active_vfcu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vfcmp & &tail | e_7_active_vfcu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vfvu <= (~_T_397 | ~(&head)) & (_T_3 & io_op_bits_active_vfconv & &tail | e_7_active_vfvu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vpu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vst & &tail | io_op_bits_active_vld &
                                                &tail) | e_7_active_vpu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vgu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vstx & &tail | io_op_bits_active_vldx &
                                                &tail | io_op_bits_active_vamo & &tail) | e_7_active_vgu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
      e_7_active_vcu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vst & &_T_0 | io_op_bits_active_vld &
                                                &_T_0 | io_op_bits_active_vstx & &_T_0 | io_op_bits_active_vldx & &_T_0 |
                                                io_op_bits_active_vamo & &_T_0) | e_7_active_vcu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21
      e_7_active_vlu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vld & &_T_1 | io_op_bits_active_vldx &
                                                &_T_1 | io_op_bits_active_vamo & &_T_2) | e_7_active_vlu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21
      e_7_active_vsu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vst & &_T_1 | io_op_bits_active_vstx &
                                                &_T_1 | io_op_bits_active_vamo & &_T_1) | e_7_active_vsu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21
      e_7_active_vqu <= (~_T_397 | ~(&head)) & (_T_3 & (io_op_bits_active_vrfirst & &tail |
                                                io_op_bits_active_vrpred & &tail | io_op_bits_active_vfdiv & &tail |
                                                io_op_bits_active_vidiv & &tail) | e_7_active_vqu);	// sequencer-master.scala:267:35, :288:26, :373:43, :389:36, :438:21, util.scala:94:11
    end
  end // always @(posedge)
  assign io_op_ready = _T;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:399:66
  assign io_master_state_valid_0 = v_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_1 = v_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_2 = v_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_3 = v_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_4 = v_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_5 = v_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_6 = v_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_valid_7 = v_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_fn_union = e_0_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_0_sreg_ss1 = e_0_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_0_sreg_ss2 = e_0_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_0_sreg_ss3 = e_0_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_0_base_vp_id = e_0_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_0_base_vp_valid = e_0_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_base_vp_scalar = e_0_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_0_base_vp_pred = e_0_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_0_base_vs1_id = e_0_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_0_base_vs1_valid = e_0_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_base_vs1_scalar = e_0_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_0_base_vs1_pred = e_0_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_0_base_vs1_prec = e_0_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_0_base_vs2_id = e_0_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_0_base_vs2_valid = e_0_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_base_vs2_scalar = e_0_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_0_base_vs2_pred = e_0_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_0_base_vs2_prec = e_0_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_0_base_vs3_id = e_0_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_0_base_vs3_valid = e_0_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_base_vs3_scalar = e_0_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_0_base_vs3_pred = e_0_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_0_base_vs3_prec = e_0_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_0_base_vd_id = e_0_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_0_base_vd_valid = e_0_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_0_base_vd_scalar = e_0_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_0_base_vd_pred = e_0_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_0_base_vd_prec = e_0_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_0_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_0_active_viu = e_0_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vipu = e_0_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vimu = e_0_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vidu = e_0_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vfmu = e_0_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vfdu = e_0_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vfcu = e_0_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vfvu = e_0_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_0_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_0_active_vpu = e_0_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vgu = e_0_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vcu = e_0_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vlu = e_0_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vsu = e_0_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_active_vqu = e_0_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_0_raw_0 = e_0_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_1 = e_0_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_2 = e_0_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_3 = e_0_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_4 = e_0_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_5 = e_0_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_6 = e_0_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_raw_7 = e_0_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_0_war_0 = e_0_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_1 = e_0_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_2 = e_0_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_3 = e_0_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_4 = e_0_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_5 = e_0_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_6 = e_0_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_war_7 = e_0_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_0_waw_0 = e_0_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_1 = e_0_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_2 = e_0_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_3 = e_0_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_4 = e_0_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_5 = e_0_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_6 = e_0_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_waw_7 = e_0_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_0_last = e_0_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_0_rports = e_0_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_0_wport_sram = e_0_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_0_wport_pred = e_0_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_1_fn_union = e_1_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_1_sreg_ss1 = e_1_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_1_sreg_ss2 = e_1_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_1_sreg_ss3 = e_1_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_1_base_vp_id = e_1_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_1_base_vp_valid = e_1_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_1_base_vp_scalar = e_1_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_1_base_vp_pred = e_1_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_1_base_vs1_id = e_1_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_1_base_vs1_valid = e_1_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_1_base_vs1_scalar = e_1_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_1_base_vs1_pred = e_1_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_1_base_vs1_prec = e_1_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_1_base_vs2_id = e_1_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_1_base_vs2_valid = e_1_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_1_base_vs2_scalar = e_1_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_1_base_vs2_pred = e_1_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_1_base_vs2_prec = e_1_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_1_base_vs3_id = e_1_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_1_base_vs3_valid = e_1_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_1_base_vs3_scalar = e_1_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_1_base_vs3_pred = e_1_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_1_base_vs3_prec = e_1_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_1_base_vd_id = e_1_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_1_base_vd_valid = e_1_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_1_base_vd_scalar = e_1_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_1_base_vd_pred = e_1_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_1_base_vd_prec = e_1_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_1_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_1_active_viu = e_1_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vipu = e_1_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vimu = e_1_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vidu = e_1_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vfmu = e_1_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vfdu = e_1_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vfcu = e_1_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vfvu = e_1_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_1_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_1_active_vpu = e_1_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vgu = e_1_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vcu = e_1_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vlu = e_1_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vsu = e_1_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_active_vqu = e_1_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_1_raw_0 = e_1_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_1 = e_1_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_2 = e_1_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_3 = e_1_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_4 = e_1_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_5 = e_1_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_6 = e_1_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_raw_7 = e_1_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_1_war_0 = e_1_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_1 = e_1_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_2 = e_1_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_3 = e_1_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_4 = e_1_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_5 = e_1_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_6 = e_1_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_war_7 = e_1_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_1_waw_0 = e_1_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_1 = e_1_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_2 = e_1_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_3 = e_1_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_4 = e_1_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_5 = e_1_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_6 = e_1_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_waw_7 = e_1_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_1_last = e_1_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_1_rports = e_1_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_1_wport_sram = e_1_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_1_wport_pred = e_1_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_2_fn_union = e_2_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_2_sreg_ss1 = e_2_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_2_sreg_ss2 = e_2_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_2_sreg_ss3 = e_2_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_2_base_vp_id = e_2_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_2_base_vp_valid = e_2_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_2_base_vp_scalar = e_2_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_2_base_vp_pred = e_2_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_2_base_vs1_id = e_2_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_2_base_vs1_valid = e_2_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_2_base_vs1_scalar = e_2_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_2_base_vs1_pred = e_2_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_2_base_vs1_prec = e_2_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_2_base_vs2_id = e_2_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_2_base_vs2_valid = e_2_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_2_base_vs2_scalar = e_2_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_2_base_vs2_pred = e_2_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_2_base_vs2_prec = e_2_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_2_base_vs3_id = e_2_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_2_base_vs3_valid = e_2_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_2_base_vs3_scalar = e_2_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_2_base_vs3_pred = e_2_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_2_base_vs3_prec = e_2_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_2_base_vd_id = e_2_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_2_base_vd_valid = e_2_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_2_base_vd_scalar = e_2_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_2_base_vd_pred = e_2_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_2_base_vd_prec = e_2_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_2_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_2_active_viu = e_2_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vipu = e_2_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vimu = e_2_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vidu = e_2_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vfmu = e_2_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vfdu = e_2_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vfcu = e_2_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vfvu = e_2_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_2_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_2_active_vpu = e_2_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vgu = e_2_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vcu = e_2_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vlu = e_2_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vsu = e_2_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_active_vqu = e_2_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_2_raw_0 = e_2_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_1 = e_2_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_2 = e_2_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_3 = e_2_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_4 = e_2_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_5 = e_2_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_6 = e_2_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_raw_7 = e_2_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_2_war_0 = e_2_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_1 = e_2_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_2 = e_2_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_3 = e_2_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_4 = e_2_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_5 = e_2_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_6 = e_2_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_war_7 = e_2_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_2_waw_0 = e_2_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_1 = e_2_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_2 = e_2_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_3 = e_2_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_4 = e_2_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_5 = e_2_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_6 = e_2_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_waw_7 = e_2_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_2_last = e_2_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_2_rports = e_2_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_2_wport_sram = e_2_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_2_wport_pred = e_2_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_3_fn_union = e_3_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_3_sreg_ss1 = e_3_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_3_sreg_ss2 = e_3_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_3_sreg_ss3 = e_3_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_3_base_vp_id = e_3_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_3_base_vp_valid = e_3_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_3_base_vp_scalar = e_3_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_3_base_vp_pred = e_3_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_3_base_vs1_id = e_3_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_3_base_vs1_valid = e_3_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_3_base_vs1_scalar = e_3_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_3_base_vs1_pred = e_3_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_3_base_vs1_prec = e_3_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_3_base_vs2_id = e_3_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_3_base_vs2_valid = e_3_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_3_base_vs2_scalar = e_3_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_3_base_vs2_pred = e_3_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_3_base_vs2_prec = e_3_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_3_base_vs3_id = e_3_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_3_base_vs3_valid = e_3_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_3_base_vs3_scalar = e_3_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_3_base_vs3_pred = e_3_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_3_base_vs3_prec = e_3_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_3_base_vd_id = e_3_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_3_base_vd_valid = e_3_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_3_base_vd_scalar = e_3_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_3_base_vd_pred = e_3_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_3_base_vd_prec = e_3_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_3_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_3_active_viu = e_3_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vipu = e_3_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vimu = e_3_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vidu = e_3_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vfmu = e_3_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vfdu = e_3_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vfcu = e_3_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vfvu = e_3_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_3_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_3_active_vpu = e_3_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vgu = e_3_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vcu = e_3_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vlu = e_3_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vsu = e_3_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_active_vqu = e_3_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_3_raw_0 = e_3_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_1 = e_3_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_2 = e_3_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_3 = e_3_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_4 = e_3_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_5 = e_3_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_6 = e_3_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_raw_7 = e_3_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_3_war_0 = e_3_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_1 = e_3_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_2 = e_3_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_3 = e_3_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_4 = e_3_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_5 = e_3_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_6 = e_3_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_war_7 = e_3_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_3_waw_0 = e_3_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_1 = e_3_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_2 = e_3_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_3 = e_3_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_4 = e_3_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_5 = e_3_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_6 = e_3_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_waw_7 = e_3_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_3_last = e_3_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_3_rports = e_3_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_3_wport_sram = e_3_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_3_wport_pred = e_3_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_4_fn_union = e_4_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_4_sreg_ss1 = e_4_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_4_sreg_ss2 = e_4_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_4_sreg_ss3 = e_4_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_4_base_vp_id = e_4_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_4_base_vp_valid = e_4_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_4_base_vp_scalar = e_4_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_4_base_vp_pred = e_4_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_4_base_vs1_id = e_4_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_4_base_vs1_valid = e_4_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_4_base_vs1_scalar = e_4_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_4_base_vs1_pred = e_4_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_4_base_vs1_prec = e_4_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_4_base_vs2_id = e_4_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_4_base_vs2_valid = e_4_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_4_base_vs2_scalar = e_4_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_4_base_vs2_pred = e_4_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_4_base_vs2_prec = e_4_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_4_base_vs3_id = e_4_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_4_base_vs3_valid = e_4_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_4_base_vs3_scalar = e_4_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_4_base_vs3_pred = e_4_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_4_base_vs3_prec = e_4_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_4_base_vd_id = e_4_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_4_base_vd_valid = e_4_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_4_base_vd_scalar = e_4_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_4_base_vd_pred = e_4_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_4_base_vd_prec = e_4_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_4_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_4_active_viu = e_4_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vipu = e_4_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vimu = e_4_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vidu = e_4_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vfmu = e_4_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vfdu = e_4_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vfcu = e_4_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vfvu = e_4_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_4_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_4_active_vpu = e_4_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vgu = e_4_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vcu = e_4_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vlu = e_4_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vsu = e_4_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_active_vqu = e_4_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_4_raw_0 = e_4_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_1 = e_4_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_2 = e_4_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_3 = e_4_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_4 = e_4_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_5 = e_4_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_6 = e_4_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_raw_7 = e_4_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_4_war_0 = e_4_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_1 = e_4_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_2 = e_4_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_3 = e_4_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_4 = e_4_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_5 = e_4_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_6 = e_4_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_war_7 = e_4_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_4_waw_0 = e_4_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_1 = e_4_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_2 = e_4_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_3 = e_4_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_4 = e_4_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_5 = e_4_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_6 = e_4_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_waw_7 = e_4_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_4_last = e_4_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_4_rports = e_4_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_4_wport_sram = e_4_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_4_wport_pred = e_4_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_5_fn_union = e_5_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_5_sreg_ss1 = e_5_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_5_sreg_ss2 = e_5_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_5_sreg_ss3 = e_5_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_5_base_vp_id = e_5_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_5_base_vp_valid = e_5_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_5_base_vp_scalar = e_5_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_5_base_vp_pred = e_5_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_5_base_vs1_id = e_5_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_5_base_vs1_valid = e_5_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_5_base_vs1_scalar = e_5_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_5_base_vs1_pred = e_5_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_5_base_vs1_prec = e_5_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_5_base_vs2_id = e_5_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_5_base_vs2_valid = e_5_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_5_base_vs2_scalar = e_5_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_5_base_vs2_pred = e_5_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_5_base_vs2_prec = e_5_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_5_base_vs3_id = e_5_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_5_base_vs3_valid = e_5_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_5_base_vs3_scalar = e_5_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_5_base_vs3_pred = e_5_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_5_base_vs3_prec = e_5_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_5_base_vd_id = e_5_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_5_base_vd_valid = e_5_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_5_base_vd_scalar = e_5_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_5_base_vd_pred = e_5_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_5_base_vd_prec = e_5_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_5_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_5_active_viu = e_5_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vipu = e_5_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vimu = e_5_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vidu = e_5_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vfmu = e_5_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vfdu = e_5_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vfcu = e_5_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vfvu = e_5_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_5_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_5_active_vpu = e_5_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vgu = e_5_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vcu = e_5_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vlu = e_5_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vsu = e_5_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_active_vqu = e_5_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_5_raw_0 = e_5_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_1 = e_5_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_2 = e_5_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_3 = e_5_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_4 = e_5_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_5 = e_5_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_6 = e_5_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_raw_7 = e_5_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_5_war_0 = e_5_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_1 = e_5_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_2 = e_5_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_3 = e_5_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_4 = e_5_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_5 = e_5_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_6 = e_5_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_war_7 = e_5_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_5_waw_0 = e_5_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_1 = e_5_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_2 = e_5_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_3 = e_5_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_4 = e_5_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_5 = e_5_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_6 = e_5_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_waw_7 = e_5_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_5_last = e_5_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_5_rports = e_5_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_5_wport_sram = e_5_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_5_wport_pred = e_5_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_6_fn_union = e_6_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_6_sreg_ss1 = e_6_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_6_sreg_ss2 = e_6_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_6_sreg_ss3 = e_6_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_6_base_vp_id = e_6_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_6_base_vp_valid = e_6_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_6_base_vp_scalar = e_6_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_6_base_vp_pred = e_6_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_6_base_vs1_id = e_6_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_6_base_vs1_valid = e_6_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_6_base_vs1_scalar = e_6_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_6_base_vs1_pred = e_6_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_6_base_vs1_prec = e_6_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_6_base_vs2_id = e_6_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_6_base_vs2_valid = e_6_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_6_base_vs2_scalar = e_6_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_6_base_vs2_pred = e_6_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_6_base_vs2_prec = e_6_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_6_base_vs3_id = e_6_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_6_base_vs3_valid = e_6_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_6_base_vs3_scalar = e_6_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_6_base_vs3_pred = e_6_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_6_base_vs3_prec = e_6_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_6_base_vd_id = e_6_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_6_base_vd_valid = e_6_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_6_base_vd_scalar = e_6_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_6_base_vd_pred = e_6_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_6_base_vd_prec = e_6_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_6_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_6_active_viu = e_6_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vipu = e_6_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vimu = e_6_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vidu = e_6_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vfmu = e_6_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vfdu = e_6_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vfcu = e_6_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vfvu = e_6_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_6_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_6_active_vpu = e_6_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vgu = e_6_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vcu = e_6_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vlu = e_6_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vsu = e_6_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_active_vqu = e_6_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_6_raw_0 = e_6_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_1 = e_6_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_2 = e_6_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_3 = e_6_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_4 = e_6_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_5 = e_6_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_6 = e_6_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_raw_7 = e_6_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_6_war_0 = e_6_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_1 = e_6_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_2 = e_6_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_3 = e_6_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_4 = e_6_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_5 = e_6_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_6 = e_6_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_war_7 = e_6_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_6_waw_0 = e_6_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_1 = e_6_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_2 = e_6_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_3 = e_6_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_4 = e_6_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_5 = e_6_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_6 = e_6_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_waw_7 = e_6_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_6_last = e_6_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_6_rports = e_6_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_6_wport_sram = e_6_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_6_wport_pred = e_6_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_e_7_fn_union = e_7_fn_union;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:289:23
  assign io_master_state_e_7_sreg_ss1 = e_7_sreg_ss1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_7_sreg_ss2 = e_7_sreg_ss2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_7_sreg_ss3 = e_7_sreg_ss3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:332:31
  assign io_master_state_e_7_base_vp_id = e_7_base_vp_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_7_base_vp_valid = e_7_base_vp_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_7_base_vp_scalar = e_7_base_vp_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_7_base_vp_pred = e_7_base_vp_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_7_base_vs1_id = e_7_base_vs1_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_7_base_vs1_valid = e_7_base_vs1_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_7_base_vs1_scalar = e_7_base_vs1_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_7_base_vs1_pred = e_7_base_vs1_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_7_base_vs1_prec = e_7_base_vs1_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_7_base_vs2_id = e_7_base_vs2_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_7_base_vs2_valid = e_7_base_vs2_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_7_base_vs2_scalar = e_7_base_vs2_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_7_base_vs2_pred = e_7_base_vs2_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_7_base_vs2_prec = e_7_base_vs2_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_7_base_vs3_id = e_7_base_vs3_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_7_base_vs3_valid = e_7_base_vs3_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_7_base_vs3_scalar = e_7_base_vs3_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_7_base_vs3_pred = e_7_base_vs3_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_7_base_vs3_prec = e_7_base_vs3_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:329:29
  assign io_master_state_e_7_base_vd_id = e_7_base_vd_id;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:141:29
  assign io_master_state_e_7_base_vd_valid = e_7_base_vd_valid;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44
  assign io_master_state_e_7_base_vd_scalar = e_7_base_vd_scalar;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:37
  assign io_master_state_e_7_base_vd_pred = e_7_base_vd_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, types-vxu.scala:119:31
  assign io_master_state_e_7_base_vd_prec = e_7_base_vd_prec;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:363:24
  assign io_master_state_e_7_rate = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_7_active_viu = e_7_active_viu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vipu = e_7_active_vipu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vimu = e_7_active_vimu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vidu = e_7_active_vidu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vfmu = e_7_active_vfmu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vfdu = e_7_active_vfdu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vfcu = e_7_active_vfcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vfvu = e_7_active_vfvu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vrpu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_7_active_vrfu = 1'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, compatibility.scala:120:12
  assign io_master_state_e_7_active_vpu = e_7_active_vpu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vgu = e_7_active_vgu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vcu = e_7_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vlu = e_7_active_vlu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vsu = e_7_active_vsu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_active_vqu = e_7_active_vqu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:288:26
  assign io_master_state_e_7_raw_0 = e_7_raw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_1 = e_7_raw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_2 = e_7_raw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_3 = e_7_raw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_4 = e_7_raw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_5 = e_7_raw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_6 = e_7_raw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_raw_7 = e_7_raw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:183:52
  assign io_master_state_e_7_war_0 = e_7_war_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_1 = e_7_war_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_2 = e_7_war_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_3 = e_7_war_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_4 = e_7_war_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_5 = e_7_war_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_6 = e_7_war_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_war_7 = e_7_war_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:184:52
  assign io_master_state_e_7_waw_0 = e_7_waw_0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_1 = e_7_waw_1;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_2 = e_7_waw_2;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_3 = e_7_waw_3;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_4 = e_7_waw_4;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_5 = e_7_waw_5;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_6 = e_7_waw_6;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_waw_7 = e_7_waw_7;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:185:52
  assign io_master_state_e_7_last = e_7_last;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:283:19
  assign io_master_state_e_7_rports = e_7_rports;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:230:21
  assign io_master_state_e_7_wport_sram = e_7_wport_sram;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:231:25
  assign io_master_state_e_7_wport_pred = e_7_wport_pred;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:232:25
  assign io_master_state_head = head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:389:36
  assign io_master_update_valid_0 = _T_385;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_1 = _T_386;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_2 = _T_387;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_3 = _T_388;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_4 = _T_389;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_5 = _T_390;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_6 = _T_391;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_valid_7 = _T_392;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_master_update_reg_0_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_291 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_4 | _T_369 ? io_op_bits_reg_vp_id : _T_361) : _T_370) :
                _T_370) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_0_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_291 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_4 | _T_345 ? io_op_bits_reg_vs2_id : _T_306) : _T_346) :
                _T_346) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_0_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_4 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_4 | _T_163 ?
                io_op_bits_reg_vs2_id : _T_124) : _T_163 ? io_op_bits_reg_vs2_id : _T_124) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_0_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_4 | _T_59 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_59 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_0_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_291 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_291 | _T_321 ? io_op_bits_reg_vd_id
                : _T_243) : _T_321 ? io_op_bits_reg_vd_id : _T_243) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_1_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_292 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_5 | _T_371 ? io_op_bits_reg_vp_id : _T_362) : _T_372) :
                _T_372) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_1_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_292 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_5 | _T_347 ? io_op_bits_reg_vs2_id : _T_307) : _T_348) :
                _T_348) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_1_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_5 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_5 | _T_164 ?
                io_op_bits_reg_vs2_id : _T_125) : _T_164 ? io_op_bits_reg_vs2_id : _T_125) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_1_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_5 | _T_60 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_60 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_1_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_292 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_292 | _T_322 ? io_op_bits_reg_vd_id
                : _T_244) : _T_322 ? io_op_bits_reg_vd_id : _T_244) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_2_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_293 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_6 | _T_373 ? io_op_bits_reg_vp_id : _T_363) : _T_374) :
                _T_374) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_2_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_293 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_6 | _T_349 ? io_op_bits_reg_vs2_id : _T_308) : _T_350) :
                _T_350) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_2_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_6 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_6 | _T_165 ?
                io_op_bits_reg_vs2_id : _T_126) : _T_165 ? io_op_bits_reg_vs2_id : _T_126) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_2_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_6 | _T_61 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_61 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_2_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_293 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_293 | _T_323 ? io_op_bits_reg_vd_id
                : _T_245) : _T_323 ? io_op_bits_reg_vd_id : _T_245) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_3_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_294 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_7 | _T_375 ? io_op_bits_reg_vp_id : _T_364) : _T_376) :
                _T_376) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_3_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_294 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_7 | _T_351 ? io_op_bits_reg_vs2_id : _T_309) : _T_352) :
                _T_352) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_3_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_7 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_7 | _T_166 ?
                io_op_bits_reg_vs2_id : _T_127) : _T_166 ? io_op_bits_reg_vs2_id : _T_127) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_3_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_7 | _T_62 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_62 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_3_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_294 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_294 | _T_324 ? io_op_bits_reg_vd_id
                : _T_246) : _T_324 ? io_op_bits_reg_vd_id : _T_246) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_4_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_295 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_8 | _T_377 ? io_op_bits_reg_vp_id : _T_365) : _T_378) :
                _T_378) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_4_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_295 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_8 | _T_353 ? io_op_bits_reg_vs2_id : _T_310) : _T_354) :
                _T_354) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_4_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_8 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_8 | _T_167 ?
                io_op_bits_reg_vs2_id : _T_128) : _T_167 ? io_op_bits_reg_vs2_id : _T_128) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_4_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_8 | _T_63 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_63 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_4_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_295 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_295 | _T_325 ? io_op_bits_reg_vd_id
                : _T_247) : _T_325 ? io_op_bits_reg_vd_id : _T_247) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_5_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_296 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_9 | _T_379 ? io_op_bits_reg_vp_id : _T_366) : _T_380) :
                _T_380) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_5_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_296 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_9 | _T_355 ? io_op_bits_reg_vs2_id : _T_311) : _T_356) :
                _T_356) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_5_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_9 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_9 | _T_168 ?
                io_op_bits_reg_vs2_id : _T_129) : _T_168 ? io_op_bits_reg_vs2_id : _T_129) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_5_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_9 | _T_64 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_64 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_5_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_296 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_296 | _T_326 ? io_op_bits_reg_vd_id
                : _T_248) : _T_326 ? io_op_bits_reg_vd_id : _T_248) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_6_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (_T_297 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (_T_10 | _T_381 ? io_op_bits_reg_vp_id : _T_367) : _T_382) :
                _T_382) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:322:41, :411:70
  assign io_master_update_reg_6_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & _T_297 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (_T_10 | _T_357 ? io_op_bits_reg_vs2_id : _T_312) : _T_358) :
                _T_358) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :356:42, :411:70
  assign io_master_update_reg_6_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & _T_10 ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (_T_10 | _T_169 ?
                io_op_bits_reg_vs2_id : _T_130) : _T_169 ? io_op_bits_reg_vs2_id : _T_130) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_6_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (_T_10 | _T_65 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_65 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:330:47, :411:70
  assign io_master_update_reg_6_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & _T_297 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (_T_297 | _T_327 ? io_op_bits_reg_vd_id
                : _T_249) : _T_327 ? io_op_bits_reg_vd_id : _T_249) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:364:41, :411:70
  assign io_master_update_reg_7_vp_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vp_valid ? (&_T_1 ? io_op_bits_reg_vp_id :
                io_op_bits_base_vp_valid ? (&tail | _T_383 ? io_op_bits_reg_vp_id : _T_368) : _T_384) :
                _T_384) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:267:35, :322:41, :411:70, util.scala:94:11
  assign io_master_update_reg_7_vs1_id = _T_3 ? (io_op_bits_active_vst & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vstx ? (io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_reg_vd_id :
                io_op_bits_base_vs2_valid ? (&tail | _T_359 ? io_op_bits_reg_vs2_id : _T_313) : _T_360) :
                _T_360) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:267:35, :330:47, :356:42, :411:70, util.scala:94:11
  assign io_master_update_reg_7_vs2_id = _T_3 ? (io_op_bits_active_vfcmp & io_op_bits_base_vs2_valid & &tail ? io_op_bits_reg_vs2_id
                : io_op_bits_active_vfdiv & io_op_bits_base_vs2_valid ? (&tail | _T_170 ?
                io_op_bits_reg_vs2_id : _T_131) : _T_170 ? io_op_bits_reg_vs2_id : _T_131) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:267:35, :330:47, :411:70, util.scala:94:11
  assign io_master_update_reg_7_vs3_id = _T_3 ? (io_op_bits_active_vfma & io_op_bits_base_vs3_valid ? (&tail | _T_66 ?
                io_op_bits_reg_vs3_id : 8'h0) : _T_66 ? io_op_bits_reg_vs3_id : 8'h0) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:267:35, :330:47, :411:70, util.scala:94:11
  assign io_master_update_reg_7_vd_id = _T_3 ? (io_op_bits_active_vld & io_op_bits_base_vd_valid & &_T_1 ? io_op_bits_reg_vd_id :
                io_op_bits_active_vldx & io_op_bits_base_vd_valid ? (&_T_1 | _T_328 ? io_op_bits_reg_vd_id
                : _T_250) : _T_328 ? io_op_bits_reg_vd_id : _T_250) : 8'h0;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:267:35, :364:41, :411:70
  assign io_pending_mem = v_0 & e_0_active_vcu | v_1 & e_1_active_vcu | v_2 & e_2_active_vcu | v_3 & e_3_active_vcu |
                v_4 & e_4_active_vcu | v_5 & e_5_active_vcu | v_6 & e_6_active_vcu | v_7 & e_7_active_vcu;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:136:44, :288:26, :446:59, :447:39
  assign io_pending_all = _T_399;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_vf_last = _T_2_398;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
  assign io_counters_memoryUOps = {1'h0, {1'h0, v_0 & (e_0_active_vgu | e_0_active_vcu | e_0_active_vlu | e_0_active_vsu)} +
                {1'h0, v_1 & (e_1_active_vgu | e_1_active_vcu | e_1_active_vlu | e_1_active_vsu)}} + {1'h0,
                {1'h0, v_2 & (e_2_active_vgu | e_2_active_vcu | e_2_active_vlu | e_2_active_vsu)} + {1'h0,
                v_3 & (e_3_active_vgu | e_3_active_vcu | e_3_active_vlu | e_3_active_vsu)}} + {1'h0, {1'h0,
                v_4 & (e_4_active_vgu | e_4_active_vcu | e_4_active_vlu | e_4_active_vsu)} + {1'h0, v_5 &
                (e_5_active_vgu | e_5_active_vcu | e_5_active_vlu | e_5_active_vsu)}} + {1'h0, {1'h0, v_6 &
                (e_6_active_vgu | e_6_active_vcu | e_6_active_vlu | e_6_active_vsu)} + {1'h0, v_7 &
                (e_7_active_vgu | e_7_active_vcu | e_7_active_vlu | e_7_active_vsu)}};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, Bitwise.scala:48:55, compatibility.scala:120:12, sequencer-master.scala:136:44, :288:26, :451:34, :452:57
  assign io_counters_arithUOps = {1'h0, {1'h0, v_0 & (e_0_active_viu | e_0_active_vimu | e_0_active_vidu | e_0_active_vfmu |
                e_0_active_vfdu | e_0_active_vfcu | e_0_active_vfvu | e_0_active_vqu)} + {1'h0, v_1 &
                (e_1_active_viu | e_1_active_vimu | e_1_active_vidu | e_1_active_vfmu | e_1_active_vfdu |
                e_1_active_vfcu | e_1_active_vfvu | e_1_active_vqu)}} + {1'h0, {1'h0, v_2 & (e_2_active_viu
                | e_2_active_vimu | e_2_active_vidu | e_2_active_vfmu | e_2_active_vfdu | e_2_active_vfcu |
                e_2_active_vfvu | e_2_active_vqu)} + {1'h0, v_3 & (e_3_active_viu | e_3_active_vimu |
                e_3_active_vidu | e_3_active_vfmu | e_3_active_vfdu | e_3_active_vfcu | e_3_active_vfvu |
                e_3_active_vqu)}} + {1'h0, {1'h0, v_4 & (e_4_active_viu | e_4_active_vimu | e_4_active_vidu
                | e_4_active_vfmu | e_4_active_vfdu | e_4_active_vfcu | e_4_active_vfvu | e_4_active_vqu)}
                + {1'h0, v_5 & (e_5_active_viu | e_5_active_vimu | e_5_active_vidu | e_5_active_vfmu |
                e_5_active_vfdu | e_5_active_vfcu | e_5_active_vfvu | e_5_active_vqu)}} + {1'h0, {1'h0, v_6
                & (e_6_active_viu | e_6_active_vimu | e_6_active_vidu | e_6_active_vfmu | e_6_active_vfdu |
                e_6_active_vfcu | e_6_active_vfvu | e_6_active_vqu)} + {1'h0, v_7 & (e_7_active_viu |
                e_7_active_vimu | e_7_active_vidu | e_7_active_vfmu | e_7_active_vfdu | e_7_active_vfcu |
                e_7_active_vfvu | e_7_active_vqu)}};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, Bitwise.scala:48:55, compatibility.scala:120:12, sequencer-master.scala:136:44, :288:26, :455:34, :457:76
  assign io_counters_predUOps = {1'h0, {1'h0, v_0 & (e_0_active_vpu | e_0_active_vipu)} + {1'h0, v_1 & (e_1_active_vpu |
                e_1_active_vipu)}} + {1'h0, {1'h0, v_2 & (e_2_active_vpu | e_2_active_vipu)} + {1'h0, v_3 &
                (e_3_active_vpu | e_3_active_vipu)}} + {1'h0, {1'h0, v_4 & (e_4_active_vpu |
                e_4_active_vipu)} + {1'h0, v_5 & (e_5_active_vpu | e_5_active_vipu)}} + {1'h0, {1'h0, v_6 &
                (e_6_active_vpu | e_6_active_vipu)} + {1'h0, v_7 & (e_7_active_vpu | e_7_active_vipu)}};	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, Bitwise.scala:48:55, compatibility.scala:120:12, sequencer-master.scala:136:44, :288:26, :461:34, :462:25
  assign io_debug_head = head;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:389:36
  assign io_debug_tail = tail;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, util.scala:94:11
  assign io_debug_maybe_full = maybe_full;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10, sequencer-master.scala:389:15
  assign io_debug_empty = _T_395;	// /Users/andrewy/wsp/circt/integration_test/Dialect/FIRRTL/Regress/HwachaSequencer.fir:6:10
endmodule

